/*-------------------------------------------------------------------------
 AES cryptographic module for FPGA on SASEBO-GIII
 
 File name   : chip_sasebo_giii_aes.v
 Version     : 1.0
 Created     : APR/02/2012
 Last update : APR/25/2013
 Desgined by : Toshihiro Katashita
 
 
 Copyright (C) 2012,2013 AIST
 
 By using this code, you agree to the following terms and conditions.
 
 This code is copyrighted by AIST ("us").
 
 Permission is hereby granted to copy, reproduce, redistribute or
 otherwise use this code as long as: there is no monetary profit gained
 specifically from the use or reproduction of this code, it is not sold,
 rented, traded or otherwise marketed, and this copyright notice is
 included prominently in any copy made.
 
 We shall not be liable for any damages, including without limitation
 direct, indirect, incidental, special or consequential damages arising
 from the use of this code.
 
 When you publish any results arising from the use of this code, we will
 appreciate it if you can cite our paper.
 (http://www.risec.aist.go.jp/project/sasebo/)
 -------------------------------------------------------------------------*/


/*-------------------------------------------------------------------------

	Implementation of Borrowed Time protection based on asynchronous circuitry
	Retained full surrounding IO framework from original source
	Comments pertaining to the countermeasure marked with 'BT'

	Designed for operating range: 2.5MHz < f < 40MHz
	however this may require tuning depending on place and route - see paper
	
  This file contains clock monitor (raising stop_detect alarm signal) and 
  delayed_edge generation circuitry, masked clearing circuitry can be found
  in AES_Composite_enc module within 

 -------------------------------------------------------------------------*/


//================================================ CHIP_SASEBO_GIII_AES
module CHIP_SASEBO_GIII_AES
  (// Local bus for GII
   lbus_di_a, lbus_do, lbus_wrn, lbus_rdn,
   lbus_clkn, lbus_rstn,

   // GPIO and LED
   gpio_startn, gpio_endn, gpio_exec, led,

   // Clock OSC
   osc_en_b);
   
   //------------------------------------------------
   // Local bus for GII
   input [15:0]  lbus_di_a;
   output [15:0] lbus_do;
   input         lbus_wrn, lbus_rdn;
   input         lbus_clkn, lbus_rstn;

   // GPIO and LED
   output        gpio_startn, gpio_endn, gpio_exec;
   output [9:0]  led;

   // Clock OSC
   output        osc_en_b;

   //------------------------------------------------
   // Internal clock
   wire         clk, rst;

   // Local bus
   reg [15:0]   lbus_a, lbus_di;
   
   // Block cipher
   wire [127:0] blk_kin, blk_din, blk_dout;
   wire         blk_krdy, blk_kvld, blk_drdy, blk_dvld;
   wire         blk_encdec, blk_en, blk_rstn, blk_busy;
   reg          blk_drdy_delay;


   //-------------------------------------------------------------------------
   //
   //	BT:	Set 'keep' attributes for each signal so EDA tools don't optimise
   // 		away signals on the delay chains or monitor circuit.
   //			
   //			delayed_edge, stop_detect - signals as labelled in paper
   //
   //			LUT outputs: EQUAL, EQUAL1, EQUAL2, EQUAL3, EQUAL4, CLK_IND
   //			for below corresponding LUTs:
   //			LUT6_1, LUT6_2, LUT6_3, LUT6_4, LUT6_5, LUT6_6
   //			all of which are input to LUT6_7, whose output is stop_detect
   //			
   //			Delay chain made up of Q_out, Q_out0, ..., Q_out2900
   //			these correspond to c0, c1, ..., cn in paper (Figure 4)
   //			they sit between delay elements: LUT1_inst, ... LUT1_inst2900
   //			taps on the chain fed are the inputs to the above listed LUTs
   //			
   //			Delayed edge delay chain made up of Q_out_dp0, ..., Q_out_dp999
   //			these correspond to s0, s1, ..., sm in paper (Figure 4)
   //			they sit between delay elements: LUT1_dpinst0, ... LUT1_dpinst1000
   //
   //			PRNG, clk_mux, & data_mux all built into AES_Composite_enc module
   //
   //-------------------------------------------------------------------------


  wire	stop_detect; // BT:	this won't be optimised away 

		  
	(* S = "true" *)
   (* KEEP = "true" *)
	wire delayed_edge;

	(* S = "true" *)  
	(* KEEP = "true" *)  
	wire CLK_IND;
	
	(* S = "true" *)  
	(* KEEP = "true" *)  
	wire EQUAL;
	
	(* S = "true" *)  
	(* KEEP = "true" *)  
	wire EQUAL1;
	
	(* S = "true" *)  
	(* KEEP = "true" *)  
	wire EQUAL2;
	
	(* S = "true" *)  
	(* KEEP = "true" *)  
	wire EQUAL3;

	(* S = "true" *)  
	(* KEEP = "true" *)  
	wire EQUAL4;
	
	(* S = "true" *)  
	(* KEEP = "true" *)  
	wire Q_out;
	
(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out0;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out2;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out3;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out4;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out5;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out6;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out7;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out8;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out9;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out10;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out11;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out12;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out13;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out14;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out15;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out16;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out17;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out18;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out19;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out20;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out21;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out22;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out23;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out24;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out25;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out26;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out27;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out28;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out29;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out30;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out31;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out32;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out33;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out34;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out35;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out36;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out37;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out38;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out39;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out40;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out41;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out42;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out43;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out44;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out45;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out46;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out47;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out48;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out49;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out50;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out51;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out52;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out53;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out54;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out55;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out56;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out57;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out58;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out59;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out60;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out61;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out62;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out63;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out64;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out65;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out66;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out67;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out68;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out69;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out70;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out71;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out72;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out73;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out74;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out75;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out76;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out77;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out78;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out79;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out80;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out81;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out82;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out83;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out84;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out85;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out86;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out87;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out88;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out89;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out90;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out91;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out92;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out93;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out94;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out95;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out96;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out97;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out98;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out99;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out100;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out101;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out102;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out103;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out104;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out105;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out106;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out107;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out108;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out109;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out110;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out111;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out112;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out113;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out114;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out115;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out116;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out117;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out118;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out119;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out120;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out121;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out122;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out123;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out124;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out125;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out126;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out127;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out128;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out129;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out130;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out131;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out132;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out133;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out134;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out135;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out136;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out137;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out138;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out139;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out140;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out141;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out142;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out143;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out144;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out145;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out146;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out147;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out148;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out149;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out150;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out151;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out152;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out153;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out154;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out155;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out156;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out157;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out158;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out159;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out160;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out161;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out162;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out163;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out164;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out165;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out166;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out167;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out168;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out169;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out170;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out171;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out172;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out173;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out174;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out175;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out176;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out177;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out178;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out179;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out180;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out181;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out182;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out183;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out184;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out185;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out186;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out187;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out188;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out189;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out190;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out191;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out192;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out193;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out194;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out195;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out196;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out197;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out198;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out199;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out200;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out201;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out202;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out203;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out204;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out205;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out206;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out207;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out208;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out209;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out210;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out211;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out212;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out213;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out214;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out215;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out216;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out217;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out218;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out219;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out220;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out221;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out222;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out223;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out224;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out225;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out226;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out227;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out228;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out229;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out230;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out231;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out232;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out233;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out234;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out235;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out236;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out237;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out238;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out239;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out240;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out241;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out242;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out243;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out244;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out245;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out246;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out247;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out248;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out249;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out250;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out251;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out252;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out253;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out254;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out255;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out256;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out257;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out258;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out259;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out260;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out261;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out262;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out263;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out264;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out265;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out266;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out267;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out268;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out269;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out270;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out271;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out272;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out273;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out274;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out275;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out276;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out277;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out278;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out279;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out280;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out281;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out282;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out283;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out284;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out285;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out286;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out287;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out288;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out289;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out290;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out291;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out292;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out293;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out294;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out295;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out296;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out297;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out298;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out299;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out300;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out301;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out302;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out303;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out304;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out305;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out306;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out307;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out308;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out309;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out310;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out311;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out312;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out313;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out314;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out315;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out316;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out317;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out318;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out319;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out320;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out321;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out322;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out323;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out324;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out325;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out326;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out327;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out328;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out329;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out330;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out331;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out332;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out333;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out334;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out335;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out336;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out337;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out338;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out339;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out340;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out341;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out342;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out343;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out344;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out345;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out346;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out347;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out348;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out349;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out350;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out351;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out352;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out353;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out354;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out355;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out356;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out357;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out358;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out359;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out360;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out361;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out362;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out363;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out364;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out365;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out366;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out367;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out368;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out369;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out370;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out371;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out372;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out373;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out374;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out375;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out376;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out377;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out378;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out379;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out380;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out381;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out382;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out383;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out384;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out385;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out386;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out387;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out388;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out389;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out390;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out391;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out392;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out393;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out394;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out395;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out396;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out397;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out398;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out399;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out400;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out401;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out402;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out403;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out404;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out405;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out406;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out407;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out408;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out409;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out410;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out411;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out412;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out413;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out414;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out415;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out416;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out417;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out418;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out419;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out420;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out421;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out422;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out423;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out424;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out425;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out426;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out427;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out428;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out429;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out430;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out431;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out432;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out433;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out434;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out435;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out436;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out437;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out438;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out439;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out440;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out441;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out442;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out443;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out444;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out445;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out446;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out447;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out448;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out449;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out450;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out451;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out452;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out453;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out454;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out455;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out456;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out457;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out458;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out459;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out460;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out461;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out462;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out463;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out464;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out465;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out466;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out467;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out468;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out469;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out470;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out471;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out472;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out473;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out474;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out475;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out476;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out477;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out478;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out479;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out480;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out481;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out482;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out483;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out484;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out485;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out486;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out487;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out488;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out489;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out490;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out491;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out492;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out493;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out494;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out495;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out496;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out497;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out498;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out499;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out500;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out501;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out502;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out503;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out504;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out505;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out506;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out507;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out508;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out509;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out510;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out511;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out512;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out513;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out514;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out515;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out516;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out517;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out518;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out519;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out520;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out521;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out522;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out523;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out524;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out525;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out526;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out527;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out528;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out529;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out530;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out531;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out532;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out533;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out534;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out535;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out536;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out537;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out538;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out539;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out540;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out541;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out542;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out543;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out544;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out545;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out546;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out547;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out548;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out549;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out550;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out551;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out552;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out553;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out554;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out555;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out556;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out557;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out558;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out559;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out560;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out561;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out562;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out563;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out564;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out565;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out566;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out567;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out568;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out569;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out570;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out571;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out572;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out573;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out574;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out575;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out576;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out577;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out578;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out579;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out580;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out581;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out582;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out583;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out584;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out585;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out586;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out587;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out588;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out589;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out590;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out591;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out592;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out593;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out594;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out595;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out596;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out597;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out598;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out599;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out600;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out601;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out602;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out603;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out604;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out605;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out606;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out607;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out608;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out609;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out610;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out611;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out612;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out613;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out614;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out615;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out616;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out617;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out618;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out619;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out620;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out621;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out622;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out623;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out624;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out625;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out626;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out627;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out628;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out629;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out630;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out631;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out632;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out633;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out634;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out635;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out636;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out637;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out638;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out639;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out640;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out641;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out642;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out643;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out644;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out645;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out646;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out647;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out648;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out649;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out650;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out651;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out652;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out653;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out654;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out655;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out656;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out657;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out658;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out659;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out660;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out661;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out662;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out663;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out664;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out665;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out666;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out667;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out668;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out669;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out670;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out671;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out672;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out673;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out674;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out675;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out676;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out677;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out678;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out679;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out680;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out681;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out682;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out683;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out684;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out685;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out686;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out687;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out688;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out689;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out690;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out691;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out692;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out693;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out694;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out695;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out696;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out697;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out698;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out699;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out700;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out701;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out702;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out703;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out704;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out705;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out706;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out707;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out708;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out709;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out710;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out711;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out712;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out713;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out714;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out715;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out716;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out717;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out718;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out719;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out720;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out721;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out722;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out723;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out724;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out725;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out726;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out727;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out728;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out729;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out730;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out731;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out732;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out733;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out734;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out735;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out736;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out737;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out738;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out739;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out740;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out741;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out742;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out743;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out744;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out745;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out746;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out747;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out748;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out749;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out750;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out751;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out752;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out753;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out754;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out755;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out756;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out757;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out758;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out759;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out760;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out761;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out762;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out763;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out764;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out765;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out766;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out767;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out768;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out769;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out770;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out771;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out772;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out773;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out774;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out775;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out776;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out777;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out778;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out779;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out780;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out781;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out782;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out783;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out784;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out785;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out786;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out787;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out788;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out789;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out790;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out791;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out792;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out793;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out794;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out795;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out796;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out797;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out798;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out799;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out800;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out801;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out802;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out803;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out804;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out805;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out806;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out807;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out808;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out809;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out810;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out811;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out812;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out813;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out814;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out815;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out816;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out817;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out818;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out819;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out820;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out821;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out822;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out823;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out824;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out825;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out826;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out827;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out828;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out829;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out830;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out831;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out832;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out833;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out834;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out835;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out836;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out837;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out838;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out839;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out840;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out841;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out842;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out843;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out844;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out845;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out846;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out847;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out848;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out849;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out850;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out851;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out852;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out853;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out854;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out855;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out856;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out857;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out858;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out859;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out860;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out861;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out862;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out863;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out864;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out865;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out866;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out867;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out868;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out869;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out870;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out871;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out872;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out873;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out874;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out875;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out876;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out877;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out878;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out879;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out880;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out881;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out882;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out883;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out884;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out885;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out886;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out887;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out888;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out889;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out890;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out891;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out892;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out893;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out894;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out895;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out896;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out897;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out898;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out899;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out900;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out901;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out902;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out903;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out904;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out905;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out906;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out907;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out908;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out909;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out910;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out911;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out912;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out913;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out914;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out915;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out916;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out917;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out918;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out919;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out920;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out921;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out922;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out923;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out924;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out925;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out926;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out927;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out928;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out929;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out930;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out931;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out932;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out933;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out934;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out935;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out936;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out937;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out938;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out939;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out940;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out941;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out942;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out943;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out944;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out945;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out946;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out947;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out948;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out949;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out950;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out951;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out952;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out953;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out954;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out955;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out956;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out957;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out958;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out959;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out960;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out961;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out962;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out963;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out964;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out965;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out966;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out967;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out968;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out969;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out970;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out971;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out972;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out973;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out974;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out975;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out976;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out977;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out978;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out979;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out980;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out981;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out982;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out983;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out984;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out985;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out986;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out987;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out988;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out989;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out990;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out991;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out992;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out993;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out994;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out995;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out996;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out997;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out998;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out999;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1000;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1001;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1002;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1003;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1004;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1005;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1006;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1007;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1008;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1009;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1010;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1011;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1012;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1013;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1014;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1015;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1016;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1017;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1018;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1019;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1020;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1021;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1022;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1023;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1024;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1025;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1026;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1027;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1028;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1029;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1030;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1031;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1032;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1033;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1034;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1035;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1036;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1037;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1038;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1039;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1040;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1041;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1042;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1043;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1044;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1045;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1046;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1047;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1048;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1049;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1050;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1051;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1052;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1053;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1054;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1055;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1056;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1057;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1058;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1059;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1060;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1061;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1062;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1063;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1064;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1065;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1066;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1067;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1068;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1069;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1070;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1071;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1072;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1073;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1074;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1075;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1076;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1077;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1078;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1079;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1080;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1081;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1082;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1083;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1084;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1085;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1086;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1087;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1088;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1089;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1090;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1091;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1092;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1093;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1094;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1095;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1096;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1097;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1098;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1099;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1100;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1101;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1102;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1103;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1104;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1105;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1106;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1107;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1108;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1109;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1110;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1111;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1112;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1113;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1114;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1115;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1116;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1117;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1118;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1119;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1120;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1121;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1122;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1123;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1124;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1125;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1126;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1127;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1128;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1129;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1130;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1131;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1132;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1133;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1134;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1135;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1136;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1137;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1138;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1139;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1140;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1141;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1142;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1143;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1144;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1145;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1146;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1147;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1148;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1149;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1150;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1151;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1152;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1153;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1154;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1155;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1156;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1157;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1158;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1159;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1160;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1161;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1162;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1163;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1164;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1165;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1166;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1167;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1168;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1169;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1170;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1171;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1172;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1173;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1174;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1175;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1176;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1177;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1178;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1179;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1180;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1181;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1182;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1183;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1184;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1185;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1186;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1187;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1188;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1189;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1190;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1191;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1192;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1193;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1194;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1195;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1196;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1197;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1198;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1199;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1200;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1201;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1202;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1203;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1204;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1205;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1206;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1207;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1208;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1209;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1210;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1211;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1212;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1213;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1214;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1215;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1216;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1217;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1218;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1219;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1220;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1221;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1222;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1223;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1224;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1225;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1226;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1227;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1228;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1229;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1230;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1231;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1232;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1233;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1234;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1235;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1236;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1237;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1238;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1239;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1240;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1241;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1242;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1243;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1244;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1245;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1246;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1247;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1248;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1249;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1250;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1251;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1252;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1253;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1254;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1255;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1256;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1257;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1258;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1259;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1260;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1261;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1262;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1263;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1264;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1265;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1266;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1267;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1268;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1269;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1270;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1271;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1272;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1273;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1274;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1275;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1276;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1277;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1278;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1279;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1280;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1281;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1282;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1283;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1284;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1285;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1286;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1287;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1288;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1289;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1290;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1291;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1292;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1293;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1294;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1295;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1296;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1297;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1298;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1299;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1300;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1301;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1302;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1303;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1304;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1305;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1306;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1307;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1308;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1309;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1310;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1311;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1312;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1313;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1314;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1315;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1316;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1317;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1318;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1319;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1320;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1321;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1322;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1323;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1324;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1325;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1326;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1327;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1328;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1329;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1330;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1331;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1332;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1333;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1334;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1335;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1336;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1337;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1338;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1339;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1340;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1341;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1342;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1343;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1344;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1345;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1346;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1347;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1348;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1349;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1350;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1351;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1352;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1353;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1354;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1355;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1356;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1357;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1358;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1359;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1360;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1361;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1362;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1363;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1364;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1365;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1366;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1367;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1368;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1369;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1370;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1371;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1372;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1373;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1374;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1375;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1376;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1377;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1378;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1379;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1380;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1381;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1382;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1383;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1384;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1385;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1386;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1387;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1388;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1389;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1390;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1391;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1392;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1393;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1394;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1395;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1396;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1397;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1398;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1399;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1400;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1401;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1402;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1403;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1404;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1405;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1406;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1407;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1408;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1409;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1410;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1411;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1412;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1413;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1414;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1415;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1416;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1417;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1418;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1419;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1420;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1421;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1422;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1423;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1424;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1425;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1426;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1427;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1428;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1429;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1430;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1431;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1432;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1433;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1434;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1435;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1436;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1437;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1438;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1439;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1440;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1441;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1442;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1443;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1444;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1445;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1446;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1447;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1448;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1449;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1450;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1451;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1452;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1453;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1454;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1455;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1456;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1457;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1458;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1459;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1460;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1461;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1462;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1463;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1464;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1465;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1466;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1467;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1468;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1469;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1470;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1471;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1472;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1473;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1474;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1475;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1476;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1477;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1478;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1479;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1480;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1481;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1482;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1483;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1484;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1485;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1486;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1487;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1488;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1489;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1490;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1491;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1492;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1493;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1494;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1495;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1496;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1497;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1498;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1499;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1500;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1501;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1502;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1503;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1504;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1505;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1506;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1507;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1508;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1509;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1510;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1511;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1512;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1513;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1514;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1515;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1516;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1517;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1518;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1519;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1520;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1521;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1522;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1523;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1524;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1525;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1526;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1527;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1528;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1529;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1530;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1531;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1532;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1533;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1534;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1535;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1536;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1537;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1538;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1539;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1540;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1541;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1542;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1543;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1544;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1545;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1546;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1547;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1548;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1549;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1550;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1551;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1552;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1553;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1554;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1555;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1556;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1557;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1558;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1559;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1560;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1561;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1562;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1563;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1564;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1565;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1566;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1567;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1568;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1569;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1570;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1571;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1572;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1573;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1574;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1575;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1576;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1577;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1578;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1579;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1580;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1581;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1582;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1583;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1584;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1585;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1586;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1587;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1588;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1589;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1590;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1591;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1592;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1593;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1594;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1595;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1596;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1597;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1598;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1599;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1600;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1601;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1602;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1603;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1604;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1605;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1606;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1607;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1608;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1609;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1610;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1611;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1612;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1613;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1614;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1615;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1616;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1617;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1618;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1619;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1620;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1621;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1622;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1623;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1624;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1625;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1626;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1627;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1628;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1629;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1630;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1631;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1632;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1633;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1634;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1635;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1636;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1637;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1638;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1639;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1640;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1641;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1642;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1643;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1644;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1645;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1646;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1647;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1648;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1649;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1650;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1651;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1652;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1653;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1654;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1655;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1656;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1657;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1658;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1659;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1660;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1661;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1662;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1663;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1664;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1665;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1666;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1667;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1668;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1669;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1670;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1671;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1672;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1673;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1674;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1675;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1676;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1677;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1678;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1679;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1680;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1681;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1682;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1683;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1684;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1685;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1686;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1687;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1688;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1689;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1690;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1691;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1692;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1693;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1694;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1695;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1696;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1697;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1698;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1699;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1700;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1701;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1702;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1703;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1704;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1705;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1706;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1707;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1708;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1709;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1710;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1711;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1712;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1713;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1714;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1715;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1716;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1717;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1718;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1719;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1720;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1721;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1722;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1723;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1724;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1725;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1726;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1727;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1728;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1729;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1730;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1731;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1732;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1733;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1734;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1735;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1736;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1737;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1738;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1739;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1740;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1741;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1742;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1743;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1744;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1745;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1746;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1747;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1748;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1749;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1750;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1751;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1752;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1753;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1754;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1755;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1756;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1757;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1758;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1759;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1760;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1761;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1762;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1763;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1764;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1765;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1766;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1767;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1768;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1769;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1770;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1771;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1772;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1773;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1774;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1775;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1776;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1777;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1778;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1779;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1780;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1781;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1782;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1783;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1784;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1785;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1786;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1787;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1788;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1789;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1790;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1791;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1792;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1793;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1794;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1795;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1796;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1797;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1798;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1799;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1800;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1801;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1802;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1803;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1804;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1805;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1806;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1807;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1808;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1809;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1810;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1811;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1812;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1813;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1814;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1815;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1816;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1817;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1818;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1819;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1820;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1821;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1822;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1823;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1824;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1825;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1826;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1827;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1828;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1829;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1830;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1831;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1832;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1833;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1834;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1835;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1836;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1837;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1838;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1839;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1840;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1841;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1842;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1843;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1844;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1845;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1846;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1847;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1848;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1849;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1850;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1851;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1852;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1853;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1854;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1855;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1856;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1857;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1858;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1859;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1860;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1861;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1862;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1863;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1864;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1865;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1866;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1867;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1868;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1869;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1870;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1871;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1872;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1873;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1874;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1875;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1876;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1877;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1878;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1879;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1880;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1881;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1882;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1883;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1884;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1885;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1886;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1887;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1888;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1889;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1890;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1891;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1892;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1893;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1894;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1895;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1896;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1897;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1898;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1899;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out1900;

	
(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out_dp0;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out_dp1;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out_dp2;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out_dp3;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out_dp4;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out_dp5;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out_dp6;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out_dp7;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out_dp8;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out_dp9;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out_dp10;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out_dp11;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out_dp12;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out_dp13;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out_dp14;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out_dp15;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out_dp16;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out_dp17;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out_dp18;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out_dp19;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out_dp20;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out_dp21;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out_dp22;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out_dp23;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out_dp24;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out_dp25;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out_dp26;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out_dp27;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out_dp28;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out_dp29;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out_dp30;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out_dp31;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out_dp32;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out_dp33;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out_dp34;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out_dp35;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out_dp36;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out_dp37;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out_dp38;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out_dp39;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out_dp40;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out_dp41;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out_dp42;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out_dp43;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out_dp44;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out_dp45;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out_dp46;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out_dp47;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out_dp48;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out_dp49;

(* S = "true" *)
	(* KEEP = "true" *)
 	wire Q_out_dp50;


    
   //------------------------------------------------
   assign led[0] = rst;
   assign led[1] = stop_detect;
   assign led[2] = 1'b0;
   assign led[3] = blk_rstn;
   assign led[4] = blk_encdec;
   assign led[5] = blk_krdy;
   assign led[6] = blk_kvld;
   assign led[7] = 1'b0;
   assign led[8] = blk_dvld;
   assign led[9] = blk_busy;

   assign osc_en_b = 1'b0;
   //------------------------------------------------
   always @(posedge clk) if (lbus_wrn)  lbus_a  <= lbus_di_a;
   always @(posedge clk) if (~lbus_wrn) lbus_di <= lbus_di_a;

   LBUS_IF lbus_if
     (.lbus_a(lbus_a), .lbus_di(lbus_di), .lbus_do(lbus_do),
      .lbus_wr(lbus_wrn), .lbus_rd(lbus_rdn),
      .blk_kin(blk_kin), .blk_din(blk_din), .blk_dout(blk_dout),
      .blk_krdy(blk_krdy), .blk_drdy(blk_drdy), 
      .blk_kvld(blk_kvld), .blk_dvld(blk_dvld),
      .blk_encdec(blk_encdec), .blk_en(blk_en), .blk_rstn(blk_rstn),
      .clk(clk), .rst(rst));

	LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst (
		.O(Q_out), // LUT general output
		.I0(clk) // LUT input
	);

	LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1 (
		.O(Q_out1), // LUT general output
		.I0(Q_out) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst2(
		.O(Q_out2), // LUT general output
		.I0(Q_out1) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst3(
		.O(Q_out3), // LUT general output
		.I0(Q_out2) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst4(
		.O(Q_out4), // LUT general output
		.I0(Q_out3) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst5(
		.O(Q_out5), // LUT general output
		.I0(Q_out4) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst6(
		.O(Q_out6), // LUT general output
		.I0(Q_out5) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst7(
		.O(Q_out7), // LUT general output
		.I0(Q_out6) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst8(
		.O(Q_out8), // LUT general output
		.I0(Q_out7) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst9(
		.O(Q_out9), // LUT general output
		.I0(Q_out8) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst10(
		.O(Q_out10), // LUT general output
		.I0(Q_out9) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst11(
		.O(Q_out11), // LUT general output
		.I0(Q_out10) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst12(
		.O(Q_out12), // LUT general output
		.I0(Q_out11) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst13(
		.O(Q_out13), // LUT general output
		.I0(Q_out12) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst14(
		.O(Q_out14), // LUT general output
		.I0(Q_out13) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst15(
		.O(Q_out15), // LUT general output
		.I0(Q_out14) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst16(
		.O(Q_out16), // LUT general output
		.I0(Q_out15) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst17(
		.O(Q_out17), // LUT general output
		.I0(Q_out16) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst18(
		.O(Q_out18), // LUT general output
		.I0(Q_out17) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst19(
		.O(Q_out19), // LUT general output
		.I0(Q_out18) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst20(
		.O(Q_out20), // LUT general output
		.I0(Q_out19) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst21(
		.O(Q_out21), // LUT general output
		.I0(Q_out20) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst22(
		.O(Q_out22), // LUT general output
		.I0(Q_out21) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst23(
		.O(Q_out23), // LUT general output
		.I0(Q_out22) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst24(
		.O(Q_out24), // LUT general output
		.I0(Q_out23) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst25(
		.O(Q_out25), // LUT general output
		.I0(Q_out24) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst26(
		.O(Q_out26), // LUT general output
		.I0(Q_out25) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst27(
		.O(Q_out27), // LUT general output
		.I0(Q_out26) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst28(
		.O(Q_out28), // LUT general output
		.I0(Q_out27) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst29(
		.O(Q_out29), // LUT general output
		.I0(Q_out28) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst30(
		.O(Q_out30), // LUT general output
		.I0(Q_out29) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst31(
		.O(Q_out31), // LUT general output
		.I0(Q_out30) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst32(
		.O(Q_out32), // LUT general output
		.I0(Q_out31) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst33(
		.O(Q_out33), // LUT general output
		.I0(Q_out32) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst34(
		.O(Q_out34), // LUT general output
		.I0(Q_out33) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst35(
		.O(Q_out35), // LUT general output
		.I0(Q_out34) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst36(
		.O(Q_out36), // LUT general output
		.I0(Q_out35) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst37(
		.O(Q_out37), // LUT general output
		.I0(Q_out36) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst38(
		.O(Q_out38), // LUT general output
		.I0(Q_out37) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst39(
		.O(Q_out39), // LUT general output
		.I0(Q_out38) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst40(
		.O(Q_out40), // LUT general output
		.I0(Q_out39) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst41(
		.O(Q_out41), // LUT general output
		.I0(Q_out40) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst42(
		.O(Q_out42), // LUT general output
		.I0(Q_out41) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst43(
		.O(Q_out43), // LUT general output
		.I0(Q_out42) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst44(
		.O(Q_out44), // LUT general output
		.I0(Q_out43) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst45(
		.O(Q_out45), // LUT general output
		.I0(Q_out44) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst46(
		.O(Q_out46), // LUT general output
		.I0(Q_out45) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst47(
		.O(Q_out47), // LUT general output
		.I0(Q_out46) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst48(
		.O(Q_out48), // LUT general output
		.I0(Q_out47) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst49(
		.O(Q_out49), // LUT general output
		.I0(Q_out48) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst50(
		.O(Q_out50), // LUT general output
		.I0(Q_out49) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst51(
		.O(Q_out51), // LUT general output
		.I0(Q_out50) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst52(
		.O(Q_out52), // LUT general output
		.I0(Q_out51) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst53(
		.O(Q_out53), // LUT general output
		.I0(Q_out52) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst54(
		.O(Q_out54), // LUT general output
		.I0(Q_out53) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst55(
		.O(Q_out55), // LUT general output
		.I0(Q_out54) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst56(
		.O(Q_out56), // LUT general output
		.I0(Q_out55) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst57(
		.O(Q_out57), // LUT general output
		.I0(Q_out56) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst58(
		.O(Q_out58), // LUT general output
		.I0(Q_out57) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst59(
		.O(Q_out59), // LUT general output
		.I0(Q_out58) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst60(
		.O(Q_out60), // LUT general output
		.I0(Q_out59) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst61(
		.O(Q_out61), // LUT general output
		.I0(Q_out60) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst62(
		.O(Q_out62), // LUT general output
		.I0(Q_out61) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst63(
		.O(Q_out63), // LUT general output
		.I0(Q_out62) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst64(
		.O(Q_out64), // LUT general output
		.I0(Q_out63) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst65(
		.O(Q_out65), // LUT general output
		.I0(Q_out64) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst66(
		.O(Q_out66), // LUT general output
		.I0(Q_out65) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst67(
		.O(Q_out67), // LUT general output
		.I0(Q_out66) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst68(
		.O(Q_out68), // LUT general output
		.I0(Q_out67) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst69(
		.O(Q_out69), // LUT general output
		.I0(Q_out68) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst70(
		.O(Q_out70), // LUT general output
		.I0(Q_out69) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst71(
		.O(Q_out71), // LUT general output
		.I0(Q_out70) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst72(
		.O(Q_out72), // LUT general output
		.I0(Q_out71) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst73(
		.O(Q_out73), // LUT general output
		.I0(Q_out72) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst74(
		.O(Q_out74), // LUT general output
		.I0(Q_out73) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst75(
		.O(Q_out75), // LUT general output
		.I0(Q_out74) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst76(
		.O(Q_out76), // LUT general output
		.I0(Q_out75) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst77(
		.O(Q_out77), // LUT general output
		.I0(Q_out76) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst78(
		.O(Q_out78), // LUT general output
		.I0(Q_out77) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst79(
		.O(Q_out79), // LUT general output
		.I0(Q_out78) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst80(
		.O(Q_out80), // LUT general output
		.I0(Q_out79) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst81(
		.O(Q_out81), // LUT general output
		.I0(Q_out80) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst82(
		.O(Q_out82), // LUT general output
		.I0(Q_out81) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst83(
		.O(Q_out83), // LUT general output
		.I0(Q_out82) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst84(
		.O(Q_out84), // LUT general output
		.I0(Q_out83) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst85(
		.O(Q_out85), // LUT general output
		.I0(Q_out84) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst86(
		.O(Q_out86), // LUT general output
		.I0(Q_out85) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst87(
		.O(Q_out87), // LUT general output
		.I0(Q_out86) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst88(
		.O(Q_out88), // LUT general output
		.I0(Q_out87) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst89(
		.O(Q_out89), // LUT general output
		.I0(Q_out88) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst90(
		.O(Q_out90), // LUT general output
		.I0(Q_out89) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst91(
		.O(Q_out91), // LUT general output
		.I0(Q_out90) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst92(
		.O(Q_out92), // LUT general output
		.I0(Q_out91) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst93(
		.O(Q_out93), // LUT general output
		.I0(Q_out92) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst94(
		.O(Q_out94), // LUT general output
		.I0(Q_out93) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst95(
		.O(Q_out95), // LUT general output
		.I0(Q_out94) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst96(
		.O(Q_out96), // LUT general output
		.I0(Q_out95) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst97(
		.O(Q_out97), // LUT general output
		.I0(Q_out96) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst98(
		.O(Q_out98), // LUT general output
		.I0(Q_out97) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst99(
		.O(Q_out99), // LUT general output
		.I0(Q_out98) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst100(
		.O(Q_out100), // LUT general output
		.I0(Q_out99) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst101(
		.O(Q_out101), // LUT general output
		.I0(Q_out100) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst102(
		.O(Q_out102), // LUT general output
		.I0(Q_out101) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst103(
		.O(Q_out103), // LUT general output
		.I0(Q_out102) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst104(
		.O(Q_out104), // LUT general output
		.I0(Q_out103) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst105(
		.O(Q_out105), // LUT general output
		.I0(Q_out104) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst106(
		.O(Q_out106), // LUT general output
		.I0(Q_out105) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst107(
		.O(Q_out107), // LUT general output
		.I0(Q_out106) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst108(
		.O(Q_out108), // LUT general output
		.I0(Q_out107) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst109(
		.O(Q_out109), // LUT general output
		.I0(Q_out108) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst110(
		.O(Q_out110), // LUT general output
		.I0(Q_out109) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst111(
		.O(Q_out111), // LUT general output
		.I0(Q_out110) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst112(
		.O(Q_out112), // LUT general output
		.I0(Q_out111) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst113(
		.O(Q_out113), // LUT general output
		.I0(Q_out112) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst114(
		.O(Q_out114), // LUT general output
		.I0(Q_out113) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst115(
		.O(Q_out115), // LUT general output
		.I0(Q_out114) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst116(
		.O(Q_out116), // LUT general output
		.I0(Q_out115) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst117(
		.O(Q_out117), // LUT general output
		.I0(Q_out116) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst118(
		.O(Q_out118), // LUT general output
		.I0(Q_out117) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst119(
		.O(Q_out119), // LUT general output
		.I0(Q_out118) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst120(
		.O(Q_out120), // LUT general output
		.I0(Q_out119) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst121(
		.O(Q_out121), // LUT general output
		.I0(Q_out120) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst122(
		.O(Q_out122), // LUT general output
		.I0(Q_out121) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst123(
		.O(Q_out123), // LUT general output
		.I0(Q_out122) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst124(
		.O(Q_out124), // LUT general output
		.I0(Q_out123) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst125(
		.O(Q_out125), // LUT general output
		.I0(Q_out124) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst126(
		.O(Q_out126), // LUT general output
		.I0(Q_out125) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst127(
		.O(Q_out127), // LUT general output
		.I0(Q_out126) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst128(
		.O(Q_out128), // LUT general output
		.I0(Q_out127) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst129(
		.O(Q_out129), // LUT general output
		.I0(Q_out128) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst130(
		.O(Q_out130), // LUT general output
		.I0(Q_out129) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst131(
		.O(Q_out131), // LUT general output
		.I0(Q_out130) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst132(
		.O(Q_out132), // LUT general output
		.I0(Q_out131) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst133(
		.O(Q_out133), // LUT general output
		.I0(Q_out132) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst134(
		.O(Q_out134), // LUT general output
		.I0(Q_out133) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst135(
		.O(Q_out135), // LUT general output
		.I0(Q_out134) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst136(
		.O(Q_out136), // LUT general output
		.I0(Q_out135) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst137(
		.O(Q_out137), // LUT general output
		.I0(Q_out136) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst138(
		.O(Q_out138), // LUT general output
		.I0(Q_out137) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst139(
		.O(Q_out139), // LUT general output
		.I0(Q_out138) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst140(
		.O(Q_out140), // LUT general output
		.I0(Q_out139) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst141(
		.O(Q_out141), // LUT general output
		.I0(Q_out140) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst142(
		.O(Q_out142), // LUT general output
		.I0(Q_out141) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst143(
		.O(Q_out143), // LUT general output
		.I0(Q_out142) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst144(
		.O(Q_out144), // LUT general output
		.I0(Q_out143) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst145(
		.O(Q_out145), // LUT general output
		.I0(Q_out144) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst146(
		.O(Q_out146), // LUT general output
		.I0(Q_out145) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst147(
		.O(Q_out147), // LUT general output
		.I0(Q_out146) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst148(
		.O(Q_out148), // LUT general output
		.I0(Q_out147) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst149(
		.O(Q_out149), // LUT general output
		.I0(Q_out148) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst150(
		.O(Q_out150), // LUT general output
		.I0(Q_out149) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst151(
		.O(Q_out151), // LUT general output
		.I0(Q_out150) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst152(
		.O(Q_out152), // LUT general output
		.I0(Q_out151) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst153(
		.O(Q_out153), // LUT general output
		.I0(Q_out152) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst154(
		.O(Q_out154), // LUT general output
		.I0(Q_out153) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst155(
		.O(Q_out155), // LUT general output
		.I0(Q_out154) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst156(
		.O(Q_out156), // LUT general output
		.I0(Q_out155) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst157(
		.O(Q_out157), // LUT general output
		.I0(Q_out156) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst158(
		.O(Q_out158), // LUT general output
		.I0(Q_out157) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst159(
		.O(Q_out159), // LUT general output
		.I0(Q_out158) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst160(
		.O(Q_out160), // LUT general output
		.I0(Q_out159) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst161(
		.O(Q_out161), // LUT general output
		.I0(Q_out160) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst162(
		.O(Q_out162), // LUT general output
		.I0(Q_out161) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst163(
		.O(Q_out163), // LUT general output
		.I0(Q_out162) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst164(
		.O(Q_out164), // LUT general output
		.I0(Q_out163) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst165(
		.O(Q_out165), // LUT general output
		.I0(Q_out164) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst166(
		.O(Q_out166), // LUT general output
		.I0(Q_out165) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst167(
		.O(Q_out167), // LUT general output
		.I0(Q_out166) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst168(
		.O(Q_out168), // LUT general output
		.I0(Q_out167) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst169(
		.O(Q_out169), // LUT general output
		.I0(Q_out168) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst170(
		.O(Q_out170), // LUT general output
		.I0(Q_out169) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst171(
		.O(Q_out171), // LUT general output
		.I0(Q_out170) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst172(
		.O(Q_out172), // LUT general output
		.I0(Q_out171) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst173(
		.O(Q_out173), // LUT general output
		.I0(Q_out172) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst174(
		.O(Q_out174), // LUT general output
		.I0(Q_out173) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst175(
		.O(Q_out175), // LUT general output
		.I0(Q_out174) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst176(
		.O(Q_out176), // LUT general output
		.I0(Q_out175) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst177(
		.O(Q_out177), // LUT general output
		.I0(Q_out176) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst178(
		.O(Q_out178), // LUT general output
		.I0(Q_out177) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst179(
		.O(Q_out179), // LUT general output
		.I0(Q_out178) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst180(
		.O(Q_out180), // LUT general output
		.I0(Q_out179) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst181(
		.O(Q_out181), // LUT general output
		.I0(Q_out180) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst182(
		.O(Q_out182), // LUT general output
		.I0(Q_out181) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst183(
		.O(Q_out183), // LUT general output
		.I0(Q_out182) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst184(
		.O(Q_out184), // LUT general output
		.I0(Q_out183) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst185(
		.O(Q_out185), // LUT general output
		.I0(Q_out184) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst186(
		.O(Q_out186), // LUT general output
		.I0(Q_out185) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst187(
		.O(Q_out187), // LUT general output
		.I0(Q_out186) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst188(
		.O(Q_out188), // LUT general output
		.I0(Q_out187) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst189(
		.O(Q_out189), // LUT general output
		.I0(Q_out188) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst190(
		.O(Q_out190), // LUT general output
		.I0(Q_out189) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst191(
		.O(Q_out191), // LUT general output
		.I0(Q_out190) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst192(
		.O(Q_out192), // LUT general output
		.I0(Q_out191) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst193(
		.O(Q_out193), // LUT general output
		.I0(Q_out192) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst194(
		.O(Q_out194), // LUT general output
		.I0(Q_out193) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst195(
		.O(Q_out195), // LUT general output
		.I0(Q_out194) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst196(
		.O(Q_out196), // LUT general output
		.I0(Q_out195) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst197(
		.O(Q_out197), // LUT general output
		.I0(Q_out196) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst198(
		.O(Q_out198), // LUT general output
		.I0(Q_out197) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst199(
		.O(Q_out199), // LUT general output
		.I0(Q_out198) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst200(
		.O(Q_out200), // LUT general output
		.I0(Q_out199) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst201(
		.O(Q_out201), // LUT general output
		.I0(Q_out200) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst202(
		.O(Q_out202), // LUT general output
		.I0(Q_out201) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst203(
		.O(Q_out203), // LUT general output
		.I0(Q_out202) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst204(
		.O(Q_out204), // LUT general output
		.I0(Q_out203) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst205(
		.O(Q_out205), // LUT general output
		.I0(Q_out204) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst206(
		.O(Q_out206), // LUT general output
		.I0(Q_out205) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst207(
		.O(Q_out207), // LUT general output
		.I0(Q_out206) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst208(
		.O(Q_out208), // LUT general output
		.I0(Q_out207) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst209(
		.O(Q_out209), // LUT general output
		.I0(Q_out208) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst210(
		.O(Q_out210), // LUT general output
		.I0(Q_out209) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst211(
		.O(Q_out211), // LUT general output
		.I0(Q_out210) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst212(
		.O(Q_out212), // LUT general output
		.I0(Q_out211) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst213(
		.O(Q_out213), // LUT general output
		.I0(Q_out212) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst214(
		.O(Q_out214), // LUT general output
		.I0(Q_out213) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst215(
		.O(Q_out215), // LUT general output
		.I0(Q_out214) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst216(
		.O(Q_out216), // LUT general output
		.I0(Q_out215) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst217(
		.O(Q_out217), // LUT general output
		.I0(Q_out216) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst218(
		.O(Q_out218), // LUT general output
		.I0(Q_out217) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst219(
		.O(Q_out219), // LUT general output
		.I0(Q_out218) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst220(
		.O(Q_out220), // LUT general output
		.I0(Q_out219) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst221(
		.O(Q_out221), // LUT general output
		.I0(Q_out220) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst222(
		.O(Q_out222), // LUT general output
		.I0(Q_out221) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst223(
		.O(Q_out223), // LUT general output
		.I0(Q_out222) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst224(
		.O(Q_out224), // LUT general output
		.I0(Q_out223) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst225(
		.O(Q_out225), // LUT general output
		.I0(Q_out224) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst226(
		.O(Q_out226), // LUT general output
		.I0(Q_out225) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst227(
		.O(Q_out227), // LUT general output
		.I0(Q_out226) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst228(
		.O(Q_out228), // LUT general output
		.I0(Q_out227) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst229(
		.O(Q_out229), // LUT general output
		.I0(Q_out228) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst230(
		.O(Q_out230), // LUT general output
		.I0(Q_out229) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst231(
		.O(Q_out231), // LUT general output
		.I0(Q_out230) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst232(
		.O(Q_out232), // LUT general output
		.I0(Q_out231) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst233(
		.O(Q_out233), // LUT general output
		.I0(Q_out232) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst234(
		.O(Q_out234), // LUT general output
		.I0(Q_out233) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst235(
		.O(Q_out235), // LUT general output
		.I0(Q_out234) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst236(
		.O(Q_out236), // LUT general output
		.I0(Q_out235) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst237(
		.O(Q_out237), // LUT general output
		.I0(Q_out236) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst238(
		.O(Q_out238), // LUT general output
		.I0(Q_out237) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst239(
		.O(Q_out239), // LUT general output
		.I0(Q_out238) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst240(
		.O(Q_out240), // LUT general output
		.I0(Q_out239) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst241(
		.O(Q_out241), // LUT general output
		.I0(Q_out240) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst242(
		.O(Q_out242), // LUT general output
		.I0(Q_out241) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst243(
		.O(Q_out243), // LUT general output
		.I0(Q_out242) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst244(
		.O(Q_out244), // LUT general output
		.I0(Q_out243) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst245(
		.O(Q_out245), // LUT general output
		.I0(Q_out244) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst246(
		.O(Q_out246), // LUT general output
		.I0(Q_out245) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst247(
		.O(Q_out247), // LUT general output
		.I0(Q_out246) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst248(
		.O(Q_out248), // LUT general output
		.I0(Q_out247) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst249(
		.O(Q_out249), // LUT general output
		.I0(Q_out248) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst250(
		.O(Q_out250), // LUT general output
		.I0(Q_out249) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst251(
		.O(Q_out251), // LUT general output
		.I0(Q_out250) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst252(
		.O(Q_out252), // LUT general output
		.I0(Q_out251) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst253(
		.O(Q_out253), // LUT general output
		.I0(Q_out252) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst254(
		.O(Q_out254), // LUT general output
		.I0(Q_out253) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst255(
		.O(Q_out255), // LUT general output
		.I0(Q_out254) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst256(
		.O(Q_out256), // LUT general output
		.I0(Q_out255) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst257(
		.O(Q_out257), // LUT general output
		.I0(Q_out256) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst258(
		.O(Q_out258), // LUT general output
		.I0(Q_out257) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst259(
		.O(Q_out259), // LUT general output
		.I0(Q_out258) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst260(
		.O(Q_out260), // LUT general output
		.I0(Q_out259) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst261(
		.O(Q_out261), // LUT general output
		.I0(Q_out260) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst262(
		.O(Q_out262), // LUT general output
		.I0(Q_out261) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst263(
		.O(Q_out263), // LUT general output
		.I0(Q_out262) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst264(
		.O(Q_out264), // LUT general output
		.I0(Q_out263) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst265(
		.O(Q_out265), // LUT general output
		.I0(Q_out264) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst266(
		.O(Q_out266), // LUT general output
		.I0(Q_out265) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst267(
		.O(Q_out267), // LUT general output
		.I0(Q_out266) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst268(
		.O(Q_out268), // LUT general output
		.I0(Q_out267) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst269(
		.O(Q_out269), // LUT general output
		.I0(Q_out268) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst270(
		.O(Q_out270), // LUT general output
		.I0(Q_out269) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst271(
		.O(Q_out271), // LUT general output
		.I0(Q_out270) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst272(
		.O(Q_out272), // LUT general output
		.I0(Q_out271) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst273(
		.O(Q_out273), // LUT general output
		.I0(Q_out272) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst274(
		.O(Q_out274), // LUT general output
		.I0(Q_out273) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst275(
		.O(Q_out275), // LUT general output
		.I0(Q_out274) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst276(
		.O(Q_out276), // LUT general output
		.I0(Q_out275) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst277(
		.O(Q_out277), // LUT general output
		.I0(Q_out276) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst278(
		.O(Q_out278), // LUT general output
		.I0(Q_out277) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst279(
		.O(Q_out279), // LUT general output
		.I0(Q_out278) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst280(
		.O(Q_out280), // LUT general output
		.I0(Q_out279) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst281(
		.O(Q_out281), // LUT general output
		.I0(Q_out280) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst282(
		.O(Q_out282), // LUT general output
		.I0(Q_out281) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst283(
		.O(Q_out283), // LUT general output
		.I0(Q_out282) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst284(
		.O(Q_out284), // LUT general output
		.I0(Q_out283) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst285(
		.O(Q_out285), // LUT general output
		.I0(Q_out284) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst286(
		.O(Q_out286), // LUT general output
		.I0(Q_out285) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst287(
		.O(Q_out287), // LUT general output
		.I0(Q_out286) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst288(
		.O(Q_out288), // LUT general output
		.I0(Q_out287) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst289(
		.O(Q_out289), // LUT general output
		.I0(Q_out288) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst290(
		.O(Q_out290), // LUT general output
		.I0(Q_out289) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst291(
		.O(Q_out291), // LUT general output
		.I0(Q_out290) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst292(
		.O(Q_out292), // LUT general output
		.I0(Q_out291) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst293(
		.O(Q_out293), // LUT general output
		.I0(Q_out292) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst294(
		.O(Q_out294), // LUT general output
		.I0(Q_out293) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst295(
		.O(Q_out295), // LUT general output
		.I0(Q_out294) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst296(
		.O(Q_out296), // LUT general output
		.I0(Q_out295) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst297(
		.O(Q_out297), // LUT general output
		.I0(Q_out296) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst298(
		.O(Q_out298), // LUT general output
		.I0(Q_out297) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst299(
		.O(Q_out299), // LUT general output
		.I0(Q_out298) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst300(
		.O(Q_out300), // LUT general output
		.I0(Q_out299) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst301(
		.O(Q_out301), // LUT general output
		.I0(Q_out300) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst302(
		.O(Q_out302), // LUT general output
		.I0(Q_out301) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst303(
		.O(Q_out303), // LUT general output
		.I0(Q_out302) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst304(
		.O(Q_out304), // LUT general output
		.I0(Q_out303) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst305(
		.O(Q_out305), // LUT general output
		.I0(Q_out304) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst306(
		.O(Q_out306), // LUT general output
		.I0(Q_out305) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst307(
		.O(Q_out307), // LUT general output
		.I0(Q_out306) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst308(
		.O(Q_out308), // LUT general output
		.I0(Q_out307) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst309(
		.O(Q_out309), // LUT general output
		.I0(Q_out308) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst310(
		.O(Q_out310), // LUT general output
		.I0(Q_out309) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst311(
		.O(Q_out311), // LUT general output
		.I0(Q_out310) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst312(
		.O(Q_out312), // LUT general output
		.I0(Q_out311) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst313(
		.O(Q_out313), // LUT general output
		.I0(Q_out312) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst314(
		.O(Q_out314), // LUT general output
		.I0(Q_out313) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst315(
		.O(Q_out315), // LUT general output
		.I0(Q_out314) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst316(
		.O(Q_out316), // LUT general output
		.I0(Q_out315) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst317(
		.O(Q_out317), // LUT general output
		.I0(Q_out316) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst318(
		.O(Q_out318), // LUT general output
		.I0(Q_out317) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst319(
		.O(Q_out319), // LUT general output
		.I0(Q_out318) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst320(
		.O(Q_out320), // LUT general output
		.I0(Q_out319) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst321(
		.O(Q_out321), // LUT general output
		.I0(Q_out320) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst322(
		.O(Q_out322), // LUT general output
		.I0(Q_out321) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst323(
		.O(Q_out323), // LUT general output
		.I0(Q_out322) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst324(
		.O(Q_out324), // LUT general output
		.I0(Q_out323) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst325(
		.O(Q_out325), // LUT general output
		.I0(Q_out324) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst326(
		.O(Q_out326), // LUT general output
		.I0(Q_out325) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst327(
		.O(Q_out327), // LUT general output
		.I0(Q_out326) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst328(
		.O(Q_out328), // LUT general output
		.I0(Q_out327) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst329(
		.O(Q_out329), // LUT general output
		.I0(Q_out328) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst330(
		.O(Q_out330), // LUT general output
		.I0(Q_out329) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst331(
		.O(Q_out331), // LUT general output
		.I0(Q_out330) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst332(
		.O(Q_out332), // LUT general output
		.I0(Q_out331) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst333(
		.O(Q_out333), // LUT general output
		.I0(Q_out332) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst334(
		.O(Q_out334), // LUT general output
		.I0(Q_out333) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst335(
		.O(Q_out335), // LUT general output
		.I0(Q_out334) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst336(
		.O(Q_out336), // LUT general output
		.I0(Q_out335) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst337(
		.O(Q_out337), // LUT general output
		.I0(Q_out336) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst338(
		.O(Q_out338), // LUT general output
		.I0(Q_out337) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst339(
		.O(Q_out339), // LUT general output
		.I0(Q_out338) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst340(
		.O(Q_out340), // LUT general output
		.I0(Q_out339) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst341(
		.O(Q_out341), // LUT general output
		.I0(Q_out340) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst342(
		.O(Q_out342), // LUT general output
		.I0(Q_out341) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst343(
		.O(Q_out343), // LUT general output
		.I0(Q_out342) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst344(
		.O(Q_out344), // LUT general output
		.I0(Q_out343) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst345(
		.O(Q_out345), // LUT general output
		.I0(Q_out344) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst346(
		.O(Q_out346), // LUT general output
		.I0(Q_out345) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst347(
		.O(Q_out347), // LUT general output
		.I0(Q_out346) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst348(
		.O(Q_out348), // LUT general output
		.I0(Q_out347) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst349(
		.O(Q_out349), // LUT general output
		.I0(Q_out348) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst350(
		.O(Q_out350), // LUT general output
		.I0(Q_out349) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst351(
		.O(Q_out351), // LUT general output
		.I0(Q_out350) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst352(
		.O(Q_out352), // LUT general output
		.I0(Q_out351) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst353(
		.O(Q_out353), // LUT general output
		.I0(Q_out352) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst354(
		.O(Q_out354), // LUT general output
		.I0(Q_out353) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst355(
		.O(Q_out355), // LUT general output
		.I0(Q_out354) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst356(
		.O(Q_out356), // LUT general output
		.I0(Q_out355) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst357(
		.O(Q_out357), // LUT general output
		.I0(Q_out356) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst358(
		.O(Q_out358), // LUT general output
		.I0(Q_out357) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst359(
		.O(Q_out359), // LUT general output
		.I0(Q_out358) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst360(
		.O(Q_out360), // LUT general output
		.I0(Q_out359) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst361(
		.O(Q_out361), // LUT general output
		.I0(Q_out360) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst362(
		.O(Q_out362), // LUT general output
		.I0(Q_out361) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst363(
		.O(Q_out363), // LUT general output
		.I0(Q_out362) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst364(
		.O(Q_out364), // LUT general output
		.I0(Q_out363) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst365(
		.O(Q_out365), // LUT general output
		.I0(Q_out364) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst366(
		.O(Q_out366), // LUT general output
		.I0(Q_out365) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst367(
		.O(Q_out367), // LUT general output
		.I0(Q_out366) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst368(
		.O(Q_out368), // LUT general output
		.I0(Q_out367) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst369(
		.O(Q_out369), // LUT general output
		.I0(Q_out368) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst370(
		.O(Q_out370), // LUT general output
		.I0(Q_out369) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst371(
		.O(Q_out371), // LUT general output
		.I0(Q_out370) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst372(
		.O(Q_out372), // LUT general output
		.I0(Q_out371) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst373(
		.O(Q_out373), // LUT general output
		.I0(Q_out372) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst374(
		.O(Q_out374), // LUT general output
		.I0(Q_out373) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst375(
		.O(Q_out375), // LUT general output
		.I0(Q_out374) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst376(
		.O(Q_out376), // LUT general output
		.I0(Q_out375) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst377(
		.O(Q_out377), // LUT general output
		.I0(Q_out376) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst378(
		.O(Q_out378), // LUT general output
		.I0(Q_out377) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst379(
		.O(Q_out379), // LUT general output
		.I0(Q_out378) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst380(
		.O(Q_out380), // LUT general output
		.I0(Q_out379) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst381(
		.O(Q_out381), // LUT general output
		.I0(Q_out380) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst382(
		.O(Q_out382), // LUT general output
		.I0(Q_out381) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst383(
		.O(Q_out383), // LUT general output
		.I0(Q_out382) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst384(
		.O(Q_out384), // LUT general output
		.I0(Q_out383) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst385(
		.O(Q_out385), // LUT general output
		.I0(Q_out384) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst386(
		.O(Q_out386), // LUT general output
		.I0(Q_out385) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst387(
		.O(Q_out387), // LUT general output
		.I0(Q_out386) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst388(
		.O(Q_out388), // LUT general output
		.I0(Q_out387) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst389(
		.O(Q_out389), // LUT general output
		.I0(Q_out388) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst390(
		.O(Q_out390), // LUT general output
		.I0(Q_out389) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst391(
		.O(Q_out391), // LUT general output
		.I0(Q_out390) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst392(
		.O(Q_out392), // LUT general output
		.I0(Q_out391) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst393(
		.O(Q_out393), // LUT general output
		.I0(Q_out392) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst394(
		.O(Q_out394), // LUT general output
		.I0(Q_out393) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst395(
		.O(Q_out395), // LUT general output
		.I0(Q_out394) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst396(
		.O(Q_out396), // LUT general output
		.I0(Q_out395) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst397(
		.O(Q_out397), // LUT general output
		.I0(Q_out396) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst398(
		.O(Q_out398), // LUT general output
		.I0(Q_out397) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst399(
		.O(Q_out399), // LUT general output
		.I0(Q_out398) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst400(
		.O(Q_out400), // LUT general output
		.I0(Q_out399) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst401(
		.O(Q_out401), // LUT general output
		.I0(Q_out400) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst402(
		.O(Q_out402), // LUT general output
		.I0(Q_out401) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst403(
		.O(Q_out403), // LUT general output
		.I0(Q_out402) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst404(
		.O(Q_out404), // LUT general output
		.I0(Q_out403) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst405(
		.O(Q_out405), // LUT general output
		.I0(Q_out404) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst406(
		.O(Q_out406), // LUT general output
		.I0(Q_out405) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst407(
		.O(Q_out407), // LUT general output
		.I0(Q_out406) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst408(
		.O(Q_out408), // LUT general output
		.I0(Q_out407) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst409(
		.O(Q_out409), // LUT general output
		.I0(Q_out408) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst410(
		.O(Q_out410), // LUT general output
		.I0(Q_out409) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst411(
		.O(Q_out411), // LUT general output
		.I0(Q_out410) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst412(
		.O(Q_out412), // LUT general output
		.I0(Q_out411) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst413(
		.O(Q_out413), // LUT general output
		.I0(Q_out412) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst414(
		.O(Q_out414), // LUT general output
		.I0(Q_out413) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst415(
		.O(Q_out415), // LUT general output
		.I0(Q_out414) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst416(
		.O(Q_out416), // LUT general output
		.I0(Q_out415) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst417(
		.O(Q_out417), // LUT general output
		.I0(Q_out416) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst418(
		.O(Q_out418), // LUT general output
		.I0(Q_out417) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst419(
		.O(Q_out419), // LUT general output
		.I0(Q_out418) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst420(
		.O(Q_out420), // LUT general output
		.I0(Q_out419) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst421(
		.O(Q_out421), // LUT general output
		.I0(Q_out420) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst422(
		.O(Q_out422), // LUT general output
		.I0(Q_out421) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst423(
		.O(Q_out423), // LUT general output
		.I0(Q_out422) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst424(
		.O(Q_out424), // LUT general output
		.I0(Q_out423) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst425(
		.O(Q_out425), // LUT general output
		.I0(Q_out424) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst426(
		.O(Q_out426), // LUT general output
		.I0(Q_out425) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst427(
		.O(Q_out427), // LUT general output
		.I0(Q_out426) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst428(
		.O(Q_out428), // LUT general output
		.I0(Q_out427) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst429(
		.O(Q_out429), // LUT general output
		.I0(Q_out428) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst430(
		.O(Q_out430), // LUT general output
		.I0(Q_out429) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst431(
		.O(Q_out431), // LUT general output
		.I0(Q_out430) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst432(
		.O(Q_out432), // LUT general output
		.I0(Q_out431) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst433(
		.O(Q_out433), // LUT general output
		.I0(Q_out432) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst434(
		.O(Q_out434), // LUT general output
		.I0(Q_out433) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst435(
		.O(Q_out435), // LUT general output
		.I0(Q_out434) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst436(
		.O(Q_out436), // LUT general output
		.I0(Q_out435) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst437(
		.O(Q_out437), // LUT general output
		.I0(Q_out436) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst438(
		.O(Q_out438), // LUT general output
		.I0(Q_out437) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst439(
		.O(Q_out439), // LUT general output
		.I0(Q_out438) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst440(
		.O(Q_out440), // LUT general output
		.I0(Q_out439) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst441(
		.O(Q_out441), // LUT general output
		.I0(Q_out440) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst442(
		.O(Q_out442), // LUT general output
		.I0(Q_out441) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst443(
		.O(Q_out443), // LUT general output
		.I0(Q_out442) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst444(
		.O(Q_out444), // LUT general output
		.I0(Q_out443) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst445(
		.O(Q_out445), // LUT general output
		.I0(Q_out444) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst446(
		.O(Q_out446), // LUT general output
		.I0(Q_out445) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst447(
		.O(Q_out447), // LUT general output
		.I0(Q_out446) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst448(
		.O(Q_out448), // LUT general output
		.I0(Q_out447) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst449(
		.O(Q_out449), // LUT general output
		.I0(Q_out448) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst450(
		.O(Q_out450), // LUT general output
		.I0(Q_out449) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst451(
		.O(Q_out451), // LUT general output
		.I0(Q_out450) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst452(
		.O(Q_out452), // LUT general output
		.I0(Q_out451) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst453(
		.O(Q_out453), // LUT general output
		.I0(Q_out452) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst454(
		.O(Q_out454), // LUT general output
		.I0(Q_out453) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst455(
		.O(Q_out455), // LUT general output
		.I0(Q_out454) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst456(
		.O(Q_out456), // LUT general output
		.I0(Q_out455) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst457(
		.O(Q_out457), // LUT general output
		.I0(Q_out456) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst458(
		.O(Q_out458), // LUT general output
		.I0(Q_out457) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst459(
		.O(Q_out459), // LUT general output
		.I0(Q_out458) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst460(
		.O(Q_out460), // LUT general output
		.I0(Q_out459) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst461(
		.O(Q_out461), // LUT general output
		.I0(Q_out460) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst462(
		.O(Q_out462), // LUT general output
		.I0(Q_out461) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst463(
		.O(Q_out463), // LUT general output
		.I0(Q_out462) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst464(
		.O(Q_out464), // LUT general output
		.I0(Q_out463) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst465(
		.O(Q_out465), // LUT general output
		.I0(Q_out464) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst466(
		.O(Q_out466), // LUT general output
		.I0(Q_out465) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst467(
		.O(Q_out467), // LUT general output
		.I0(Q_out466) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst468(
		.O(Q_out468), // LUT general output
		.I0(Q_out467) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst469(
		.O(Q_out469), // LUT general output
		.I0(Q_out468) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst470(
		.O(Q_out470), // LUT general output
		.I0(Q_out469) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst471(
		.O(Q_out471), // LUT general output
		.I0(Q_out470) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst472(
		.O(Q_out472), // LUT general output
		.I0(Q_out471) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst473(
		.O(Q_out473), // LUT general output
		.I0(Q_out472) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst474(
		.O(Q_out474), // LUT general output
		.I0(Q_out473) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst475(
		.O(Q_out475), // LUT general output
		.I0(Q_out474) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst476(
		.O(Q_out476), // LUT general output
		.I0(Q_out475) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst477(
		.O(Q_out477), // LUT general output
		.I0(Q_out476) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst478(
		.O(Q_out478), // LUT general output
		.I0(Q_out477) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst479(
		.O(Q_out479), // LUT general output
		.I0(Q_out478) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst480(
		.O(Q_out480), // LUT general output
		.I0(Q_out479) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst481(
		.O(Q_out481), // LUT general output
		.I0(Q_out480) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst482(
		.O(Q_out482), // LUT general output
		.I0(Q_out481) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst483(
		.O(Q_out483), // LUT general output
		.I0(Q_out482) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst484(
		.O(Q_out484), // LUT general output
		.I0(Q_out483) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst485(
		.O(Q_out485), // LUT general output
		.I0(Q_out484) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst486(
		.O(Q_out486), // LUT general output
		.I0(Q_out485) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst487(
		.O(Q_out487), // LUT general output
		.I0(Q_out486) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst488(
		.O(Q_out488), // LUT general output
		.I0(Q_out487) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst489(
		.O(Q_out489), // LUT general output
		.I0(Q_out488) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst490(
		.O(Q_out490), // LUT general output
		.I0(Q_out489) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst491(
		.O(Q_out491), // LUT general output
		.I0(Q_out490) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst492(
		.O(Q_out492), // LUT general output
		.I0(Q_out491) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst493(
		.O(Q_out493), // LUT general output
		.I0(Q_out492) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst494(
		.O(Q_out494), // LUT general output
		.I0(Q_out493) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst495(
		.O(Q_out495), // LUT general output
		.I0(Q_out494) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst496(
		.O(Q_out496), // LUT general output
		.I0(Q_out495) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst497(
		.O(Q_out497), // LUT general output
		.I0(Q_out496) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst498(
		.O(Q_out498), // LUT general output
		.I0(Q_out497) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst499(
		.O(Q_out499), // LUT general output
		.I0(Q_out498) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst500(
		.O(Q_out500), // LUT general output
		.I0(Q_out499) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst501(
		.O(Q_out501), // LUT general output
		.I0(Q_out500) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst502(
		.O(Q_out502), // LUT general output
		.I0(Q_out501) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst503(
		.O(Q_out503), // LUT general output
		.I0(Q_out502) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst504(
		.O(Q_out504), // LUT general output
		.I0(Q_out503) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst505(
		.O(Q_out505), // LUT general output
		.I0(Q_out504) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst506(
		.O(Q_out506), // LUT general output
		.I0(Q_out505) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst507(
		.O(Q_out507), // LUT general output
		.I0(Q_out506) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst508(
		.O(Q_out508), // LUT general output
		.I0(Q_out507) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst509(
		.O(Q_out509), // LUT general output
		.I0(Q_out508) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst510(
		.O(Q_out510), // LUT general output
		.I0(Q_out509) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst511(
		.O(Q_out511), // LUT general output
		.I0(Q_out510) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst512(
		.O(Q_out512), // LUT general output
		.I0(Q_out511) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst513(
		.O(Q_out513), // LUT general output
		.I0(Q_out512) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst514(
		.O(Q_out514), // LUT general output
		.I0(Q_out513) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst515(
		.O(Q_out515), // LUT general output
		.I0(Q_out514) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst516(
		.O(Q_out516), // LUT general output
		.I0(Q_out515) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst517(
		.O(Q_out517), // LUT general output
		.I0(Q_out516) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst518(
		.O(Q_out518), // LUT general output
		.I0(Q_out517) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst519(
		.O(Q_out519), // LUT general output
		.I0(Q_out518) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst520(
		.O(Q_out520), // LUT general output
		.I0(Q_out519) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst521(
		.O(Q_out521), // LUT general output
		.I0(Q_out520) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst522(
		.O(Q_out522), // LUT general output
		.I0(Q_out521) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst523(
		.O(Q_out523), // LUT general output
		.I0(Q_out522) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst524(
		.O(Q_out524), // LUT general output
		.I0(Q_out523) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst525(
		.O(Q_out525), // LUT general output
		.I0(Q_out524) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst526(
		.O(Q_out526), // LUT general output
		.I0(Q_out525) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst527(
		.O(Q_out527), // LUT general output
		.I0(Q_out526) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst528(
		.O(Q_out528), // LUT general output
		.I0(Q_out527) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst529(
		.O(Q_out529), // LUT general output
		.I0(Q_out528) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst530(
		.O(Q_out530), // LUT general output
		.I0(Q_out529) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst531(
		.O(Q_out531), // LUT general output
		.I0(Q_out530) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst532(
		.O(Q_out532), // LUT general output
		.I0(Q_out531) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst533(
		.O(Q_out533), // LUT general output
		.I0(Q_out532) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst534(
		.O(Q_out534), // LUT general output
		.I0(Q_out533) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst535(
		.O(Q_out535), // LUT general output
		.I0(Q_out534) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst536(
		.O(Q_out536), // LUT general output
		.I0(Q_out535) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst537(
		.O(Q_out537), // LUT general output
		.I0(Q_out536) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst538(
		.O(Q_out538), // LUT general output
		.I0(Q_out537) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst539(
		.O(Q_out539), // LUT general output
		.I0(Q_out538) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst540(
		.O(Q_out540), // LUT general output
		.I0(Q_out539) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst541(
		.O(Q_out541), // LUT general output
		.I0(Q_out540) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst542(
		.O(Q_out542), // LUT general output
		.I0(Q_out541) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst543(
		.O(Q_out543), // LUT general output
		.I0(Q_out542) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst544(
		.O(Q_out544), // LUT general output
		.I0(Q_out543) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst545(
		.O(Q_out545), // LUT general output
		.I0(Q_out544) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst546(
		.O(Q_out546), // LUT general output
		.I0(Q_out545) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst547(
		.O(Q_out547), // LUT general output
		.I0(Q_out546) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst548(
		.O(Q_out548), // LUT general output
		.I0(Q_out547) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst549(
		.O(Q_out549), // LUT general output
		.I0(Q_out548) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst550(
		.O(Q_out550), // LUT general output
		.I0(Q_out549) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst551(
		.O(Q_out551), // LUT general output
		.I0(Q_out550) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst552(
		.O(Q_out552), // LUT general output
		.I0(Q_out551) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst553(
		.O(Q_out553), // LUT general output
		.I0(Q_out552) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst554(
		.O(Q_out554), // LUT general output
		.I0(Q_out553) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst555(
		.O(Q_out555), // LUT general output
		.I0(Q_out554) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst556(
		.O(Q_out556), // LUT general output
		.I0(Q_out555) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst557(
		.O(Q_out557), // LUT general output
		.I0(Q_out556) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst558(
		.O(Q_out558), // LUT general output
		.I0(Q_out557) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst559(
		.O(Q_out559), // LUT general output
		.I0(Q_out558) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst560(
		.O(Q_out560), // LUT general output
		.I0(Q_out559) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst561(
		.O(Q_out561), // LUT general output
		.I0(Q_out560) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst562(
		.O(Q_out562), // LUT general output
		.I0(Q_out561) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst563(
		.O(Q_out563), // LUT general output
		.I0(Q_out562) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst564(
		.O(Q_out564), // LUT general output
		.I0(Q_out563) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst565(
		.O(Q_out565), // LUT general output
		.I0(Q_out564) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst566(
		.O(Q_out566), // LUT general output
		.I0(Q_out565) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst567(
		.O(Q_out567), // LUT general output
		.I0(Q_out566) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst568(
		.O(Q_out568), // LUT general output
		.I0(Q_out567) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst569(
		.O(Q_out569), // LUT general output
		.I0(Q_out568) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst570(
		.O(Q_out570), // LUT general output
		.I0(Q_out569) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst571(
		.O(Q_out571), // LUT general output
		.I0(Q_out570) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst572(
		.O(Q_out572), // LUT general output
		.I0(Q_out571) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst573(
		.O(Q_out573), // LUT general output
		.I0(Q_out572) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst574(
		.O(Q_out574), // LUT general output
		.I0(Q_out573) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst575(
		.O(Q_out575), // LUT general output
		.I0(Q_out574) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst576(
		.O(Q_out576), // LUT general output
		.I0(Q_out575) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst577(
		.O(Q_out577), // LUT general output
		.I0(Q_out576) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst578(
		.O(Q_out578), // LUT general output
		.I0(Q_out577) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst579(
		.O(Q_out579), // LUT general output
		.I0(Q_out578) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst580(
		.O(Q_out580), // LUT general output
		.I0(Q_out579) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst581(
		.O(Q_out581), // LUT general output
		.I0(Q_out580) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst582(
		.O(Q_out582), // LUT general output
		.I0(Q_out581) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst583(
		.O(Q_out583), // LUT general output
		.I0(Q_out582) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst584(
		.O(Q_out584), // LUT general output
		.I0(Q_out583) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst585(
		.O(Q_out585), // LUT general output
		.I0(Q_out584) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst586(
		.O(Q_out586), // LUT general output
		.I0(Q_out585) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst587(
		.O(Q_out587), // LUT general output
		.I0(Q_out586) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst588(
		.O(Q_out588), // LUT general output
		.I0(Q_out587) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst589(
		.O(Q_out589), // LUT general output
		.I0(Q_out588) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst590(
		.O(Q_out590), // LUT general output
		.I0(Q_out589) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst591(
		.O(Q_out591), // LUT general output
		.I0(Q_out590) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst592(
		.O(Q_out592), // LUT general output
		.I0(Q_out591) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst593(
		.O(Q_out593), // LUT general output
		.I0(Q_out592) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst594(
		.O(Q_out594), // LUT general output
		.I0(Q_out593) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst595(
		.O(Q_out595), // LUT general output
		.I0(Q_out594) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst596(
		.O(Q_out596), // LUT general output
		.I0(Q_out595) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst597(
		.O(Q_out597), // LUT general output
		.I0(Q_out596) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst598(
		.O(Q_out598), // LUT general output
		.I0(Q_out597) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst599(
		.O(Q_out599), // LUT general output
		.I0(Q_out598) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst600(
		.O(Q_out600), // LUT general output
		.I0(Q_out599) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst601(
		.O(Q_out601), // LUT general output
		.I0(Q_out600) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst602(
		.O(Q_out602), // LUT general output
		.I0(Q_out601) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst603(
		.O(Q_out603), // LUT general output
		.I0(Q_out602) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst604(
		.O(Q_out604), // LUT general output
		.I0(Q_out603) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst605(
		.O(Q_out605), // LUT general output
		.I0(Q_out604) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst606(
		.O(Q_out606), // LUT general output
		.I0(Q_out605) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst607(
		.O(Q_out607), // LUT general output
		.I0(Q_out606) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst608(
		.O(Q_out608), // LUT general output
		.I0(Q_out607) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst609(
		.O(Q_out609), // LUT general output
		.I0(Q_out608) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst610(
		.O(Q_out610), // LUT general output
		.I0(Q_out609) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst611(
		.O(Q_out611), // LUT general output
		.I0(Q_out610) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst612(
		.O(Q_out612), // LUT general output
		.I0(Q_out611) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst613(
		.O(Q_out613), // LUT general output
		.I0(Q_out612) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst614(
		.O(Q_out614), // LUT general output
		.I0(Q_out613) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst615(
		.O(Q_out615), // LUT general output
		.I0(Q_out614) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst616(
		.O(Q_out616), // LUT general output
		.I0(Q_out615) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst617(
		.O(Q_out617), // LUT general output
		.I0(Q_out616) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst618(
		.O(Q_out618), // LUT general output
		.I0(Q_out617) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst619(
		.O(Q_out619), // LUT general output
		.I0(Q_out618) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst620(
		.O(Q_out620), // LUT general output
		.I0(Q_out619) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst621(
		.O(Q_out621), // LUT general output
		.I0(Q_out620) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst622(
		.O(Q_out622), // LUT general output
		.I0(Q_out621) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst623(
		.O(Q_out623), // LUT general output
		.I0(Q_out622) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst624(
		.O(Q_out624), // LUT general output
		.I0(Q_out623) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst625(
		.O(Q_out625), // LUT general output
		.I0(Q_out624) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst626(
		.O(Q_out626), // LUT general output
		.I0(Q_out625) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst627(
		.O(Q_out627), // LUT general output
		.I0(Q_out626) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst628(
		.O(Q_out628), // LUT general output
		.I0(Q_out627) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst629(
		.O(Q_out629), // LUT general output
		.I0(Q_out628) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst630(
		.O(Q_out630), // LUT general output
		.I0(Q_out629) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst631(
		.O(Q_out631), // LUT general output
		.I0(Q_out630) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst632(
		.O(Q_out632), // LUT general output
		.I0(Q_out631) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst633(
		.O(Q_out633), // LUT general output
		.I0(Q_out632) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst634(
		.O(Q_out634), // LUT general output
		.I0(Q_out633) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst635(
		.O(Q_out635), // LUT general output
		.I0(Q_out634) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst636(
		.O(Q_out636), // LUT general output
		.I0(Q_out635) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst637(
		.O(Q_out637), // LUT general output
		.I0(Q_out636) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst638(
		.O(Q_out638), // LUT general output
		.I0(Q_out637) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst639(
		.O(Q_out639), // LUT general output
		.I0(Q_out638) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst640(
		.O(Q_out640), // LUT general output
		.I0(Q_out639) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst641(
		.O(Q_out641), // LUT general output
		.I0(Q_out640) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst642(
		.O(Q_out642), // LUT general output
		.I0(Q_out641) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst643(
		.O(Q_out643), // LUT general output
		.I0(Q_out642) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst644(
		.O(Q_out644), // LUT general output
		.I0(Q_out643) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst645(
		.O(Q_out645), // LUT general output
		.I0(Q_out644) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst646(
		.O(Q_out646), // LUT general output
		.I0(Q_out645) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst647(
		.O(Q_out647), // LUT general output
		.I0(Q_out646) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst648(
		.O(Q_out648), // LUT general output
		.I0(Q_out647) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst649(
		.O(Q_out649), // LUT general output
		.I0(Q_out648) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst650(
		.O(Q_out650), // LUT general output
		.I0(Q_out649) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst651(
		.O(Q_out651), // LUT general output
		.I0(Q_out650) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst652(
		.O(Q_out652), // LUT general output
		.I0(Q_out651) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst653(
		.O(Q_out653), // LUT general output
		.I0(Q_out652) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst654(
		.O(Q_out654), // LUT general output
		.I0(Q_out653) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst655(
		.O(Q_out655), // LUT general output
		.I0(Q_out654) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst656(
		.O(Q_out656), // LUT general output
		.I0(Q_out655) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst657(
		.O(Q_out657), // LUT general output
		.I0(Q_out656) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst658(
		.O(Q_out658), // LUT general output
		.I0(Q_out657) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst659(
		.O(Q_out659), // LUT general output
		.I0(Q_out658) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst660(
		.O(Q_out660), // LUT general output
		.I0(Q_out659) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst661(
		.O(Q_out661), // LUT general output
		.I0(Q_out660) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst662(
		.O(Q_out662), // LUT general output
		.I0(Q_out661) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst663(
		.O(Q_out663), // LUT general output
		.I0(Q_out662) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst664(
		.O(Q_out664), // LUT general output
		.I0(Q_out663) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst665(
		.O(Q_out665), // LUT general output
		.I0(Q_out664) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst666(
		.O(Q_out666), // LUT general output
		.I0(Q_out665) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst667(
		.O(Q_out667), // LUT general output
		.I0(Q_out666) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst668(
		.O(Q_out668), // LUT general output
		.I0(Q_out667) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst669(
		.O(Q_out669), // LUT general output
		.I0(Q_out668) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst670(
		.O(Q_out670), // LUT general output
		.I0(Q_out669) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst671(
		.O(Q_out671), // LUT general output
		.I0(Q_out670) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst672(
		.O(Q_out672), // LUT general output
		.I0(Q_out671) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst673(
		.O(Q_out673), // LUT general output
		.I0(Q_out672) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst674(
		.O(Q_out674), // LUT general output
		.I0(Q_out673) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst675(
		.O(Q_out675), // LUT general output
		.I0(Q_out674) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst676(
		.O(Q_out676), // LUT general output
		.I0(Q_out675) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst677(
		.O(Q_out677), // LUT general output
		.I0(Q_out676) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst678(
		.O(Q_out678), // LUT general output
		.I0(Q_out677) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst679(
		.O(Q_out679), // LUT general output
		.I0(Q_out678) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst680(
		.O(Q_out680), // LUT general output
		.I0(Q_out679) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst681(
		.O(Q_out681), // LUT general output
		.I0(Q_out680) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst682(
		.O(Q_out682), // LUT general output
		.I0(Q_out681) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst683(
		.O(Q_out683), // LUT general output
		.I0(Q_out682) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst684(
		.O(Q_out684), // LUT general output
		.I0(Q_out683) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst685(
		.O(Q_out685), // LUT general output
		.I0(Q_out684) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst686(
		.O(Q_out686), // LUT general output
		.I0(Q_out685) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst687(
		.O(Q_out687), // LUT general output
		.I0(Q_out686) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst688(
		.O(Q_out688), // LUT general output
		.I0(Q_out687) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst689(
		.O(Q_out689), // LUT general output
		.I0(Q_out688) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst690(
		.O(Q_out690), // LUT general output
		.I0(Q_out689) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst691(
		.O(Q_out691), // LUT general output
		.I0(Q_out690) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst692(
		.O(Q_out692), // LUT general output
		.I0(Q_out691) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst693(
		.O(Q_out693), // LUT general output
		.I0(Q_out692) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst694(
		.O(Q_out694), // LUT general output
		.I0(Q_out693) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst695(
		.O(Q_out695), // LUT general output
		.I0(Q_out694) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst696(
		.O(Q_out696), // LUT general output
		.I0(Q_out695) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst697(
		.O(Q_out697), // LUT general output
		.I0(Q_out696) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst698(
		.O(Q_out698), // LUT general output
		.I0(Q_out697) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst699(
		.O(Q_out699), // LUT general output
		.I0(Q_out698) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst700(
		.O(Q_out700), // LUT general output
		.I0(Q_out699) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst701(
		.O(Q_out701), // LUT general output
		.I0(Q_out700) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst702(
		.O(Q_out702), // LUT general output
		.I0(Q_out701) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst703(
		.O(Q_out703), // LUT general output
		.I0(Q_out702) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst704(
		.O(Q_out704), // LUT general output
		.I0(Q_out703) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst705(
		.O(Q_out705), // LUT general output
		.I0(Q_out704) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst706(
		.O(Q_out706), // LUT general output
		.I0(Q_out705) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst707(
		.O(Q_out707), // LUT general output
		.I0(Q_out706) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst708(
		.O(Q_out708), // LUT general output
		.I0(Q_out707) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst709(
		.O(Q_out709), // LUT general output
		.I0(Q_out708) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst710(
		.O(Q_out710), // LUT general output
		.I0(Q_out709) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst711(
		.O(Q_out711), // LUT general output
		.I0(Q_out710) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst712(
		.O(Q_out712), // LUT general output
		.I0(Q_out711) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst713(
		.O(Q_out713), // LUT general output
		.I0(Q_out712) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst714(
		.O(Q_out714), // LUT general output
		.I0(Q_out713) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst715(
		.O(Q_out715), // LUT general output
		.I0(Q_out714) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst716(
		.O(Q_out716), // LUT general output
		.I0(Q_out715) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst717(
		.O(Q_out717), // LUT general output
		.I0(Q_out716) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst718(
		.O(Q_out718), // LUT general output
		.I0(Q_out717) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst719(
		.O(Q_out719), // LUT general output
		.I0(Q_out718) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst720(
		.O(Q_out720), // LUT general output
		.I0(Q_out719) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst721(
		.O(Q_out721), // LUT general output
		.I0(Q_out720) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst722(
		.O(Q_out722), // LUT general output
		.I0(Q_out721) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst723(
		.O(Q_out723), // LUT general output
		.I0(Q_out722) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst724(
		.O(Q_out724), // LUT general output
		.I0(Q_out723) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst725(
		.O(Q_out725), // LUT general output
		.I0(Q_out724) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst726(
		.O(Q_out726), // LUT general output
		.I0(Q_out725) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst727(
		.O(Q_out727), // LUT general output
		.I0(Q_out726) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst728(
		.O(Q_out728), // LUT general output
		.I0(Q_out727) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst729(
		.O(Q_out729), // LUT general output
		.I0(Q_out728) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst730(
		.O(Q_out730), // LUT general output
		.I0(Q_out729) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst731(
		.O(Q_out731), // LUT general output
		.I0(Q_out730) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst732(
		.O(Q_out732), // LUT general output
		.I0(Q_out731) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst733(
		.O(Q_out733), // LUT general output
		.I0(Q_out732) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst734(
		.O(Q_out734), // LUT general output
		.I0(Q_out733) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst735(
		.O(Q_out735), // LUT general output
		.I0(Q_out734) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst736(
		.O(Q_out736), // LUT general output
		.I0(Q_out735) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst737(
		.O(Q_out737), // LUT general output
		.I0(Q_out736) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst738(
		.O(Q_out738), // LUT general output
		.I0(Q_out737) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst739(
		.O(Q_out739), // LUT general output
		.I0(Q_out738) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst740(
		.O(Q_out740), // LUT general output
		.I0(Q_out739) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst741(
		.O(Q_out741), // LUT general output
		.I0(Q_out740) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst742(
		.O(Q_out742), // LUT general output
		.I0(Q_out741) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst743(
		.O(Q_out743), // LUT general output
		.I0(Q_out742) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst744(
		.O(Q_out744), // LUT general output
		.I0(Q_out743) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst745(
		.O(Q_out745), // LUT general output
		.I0(Q_out744) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst746(
		.O(Q_out746), // LUT general output
		.I0(Q_out745) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst747(
		.O(Q_out747), // LUT general output
		.I0(Q_out746) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst748(
		.O(Q_out748), // LUT general output
		.I0(Q_out747) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst749(
		.O(Q_out749), // LUT general output
		.I0(Q_out748) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst750(
		.O(Q_out750), // LUT general output
		.I0(Q_out749) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst751(
		.O(Q_out751), // LUT general output
		.I0(Q_out750) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst752(
		.O(Q_out752), // LUT general output
		.I0(Q_out751) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst753(
		.O(Q_out753), // LUT general output
		.I0(Q_out752) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst754(
		.O(Q_out754), // LUT general output
		.I0(Q_out753) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst755(
		.O(Q_out755), // LUT general output
		.I0(Q_out754) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst756(
		.O(Q_out756), // LUT general output
		.I0(Q_out755) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst757(
		.O(Q_out757), // LUT general output
		.I0(Q_out756) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst758(
		.O(Q_out758), // LUT general output
		.I0(Q_out757) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst759(
		.O(Q_out759), // LUT general output
		.I0(Q_out758) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst760(
		.O(Q_out760), // LUT general output
		.I0(Q_out759) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst761(
		.O(Q_out761), // LUT general output
		.I0(Q_out760) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst762(
		.O(Q_out762), // LUT general output
		.I0(Q_out761) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst763(
		.O(Q_out763), // LUT general output
		.I0(Q_out762) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst764(
		.O(Q_out764), // LUT general output
		.I0(Q_out763) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst765(
		.O(Q_out765), // LUT general output
		.I0(Q_out764) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst766(
		.O(Q_out766), // LUT general output
		.I0(Q_out765) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst767(
		.O(Q_out767), // LUT general output
		.I0(Q_out766) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst768(
		.O(Q_out768), // LUT general output
		.I0(Q_out767) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst769(
		.O(Q_out769), // LUT general output
		.I0(Q_out768) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst770(
		.O(Q_out770), // LUT general output
		.I0(Q_out769) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst771(
		.O(Q_out771), // LUT general output
		.I0(Q_out770) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst772(
		.O(Q_out772), // LUT general output
		.I0(Q_out771) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst773(
		.O(Q_out773), // LUT general output
		.I0(Q_out772) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst774(
		.O(Q_out774), // LUT general output
		.I0(Q_out773) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst775(
		.O(Q_out775), // LUT general output
		.I0(Q_out774) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst776(
		.O(Q_out776), // LUT general output
		.I0(Q_out775) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst777(
		.O(Q_out777), // LUT general output
		.I0(Q_out776) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst778(
		.O(Q_out778), // LUT general output
		.I0(Q_out777) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst779(
		.O(Q_out779), // LUT general output
		.I0(Q_out778) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst780(
		.O(Q_out780), // LUT general output
		.I0(Q_out779) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst781(
		.O(Q_out781), // LUT general output
		.I0(Q_out780) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst782(
		.O(Q_out782), // LUT general output
		.I0(Q_out781) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst783(
		.O(Q_out783), // LUT general output
		.I0(Q_out782) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst784(
		.O(Q_out784), // LUT general output
		.I0(Q_out783) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst785(
		.O(Q_out785), // LUT general output
		.I0(Q_out784) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst786(
		.O(Q_out786), // LUT general output
		.I0(Q_out785) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst787(
		.O(Q_out787), // LUT general output
		.I0(Q_out786) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst788(
		.O(Q_out788), // LUT general output
		.I0(Q_out787) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst789(
		.O(Q_out789), // LUT general output
		.I0(Q_out788) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst790(
		.O(Q_out790), // LUT general output
		.I0(Q_out789) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst791(
		.O(Q_out791), // LUT general output
		.I0(Q_out790) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst792(
		.O(Q_out792), // LUT general output
		.I0(Q_out791) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst793(
		.O(Q_out793), // LUT general output
		.I0(Q_out792) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst794(
		.O(Q_out794), // LUT general output
		.I0(Q_out793) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst795(
		.O(Q_out795), // LUT general output
		.I0(Q_out794) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst796(
		.O(Q_out796), // LUT general output
		.I0(Q_out795) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst797(
		.O(Q_out797), // LUT general output
		.I0(Q_out796) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst798(
		.O(Q_out798), // LUT general output
		.I0(Q_out797) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst799(
		.O(Q_out799), // LUT general output
		.I0(Q_out798) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst800(
		.O(Q_out800), // LUT general output
		.I0(Q_out799) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst801(
		.O(Q_out801), // LUT general output
		.I0(Q_out800) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst802(
		.O(Q_out802), // LUT general output
		.I0(Q_out801) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst803(
		.O(Q_out803), // LUT general output
		.I0(Q_out802) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst804(
		.O(Q_out804), // LUT general output
		.I0(Q_out803) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst805(
		.O(Q_out805), // LUT general output
		.I0(Q_out804) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst806(
		.O(Q_out806), // LUT general output
		.I0(Q_out805) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst807(
		.O(Q_out807), // LUT general output
		.I0(Q_out806) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst808(
		.O(Q_out808), // LUT general output
		.I0(Q_out807) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst809(
		.O(Q_out809), // LUT general output
		.I0(Q_out808) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst810(
		.O(Q_out810), // LUT general output
		.I0(Q_out809) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst811(
		.O(Q_out811), // LUT general output
		.I0(Q_out810) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst812(
		.O(Q_out812), // LUT general output
		.I0(Q_out811) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst813(
		.O(Q_out813), // LUT general output
		.I0(Q_out812) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst814(
		.O(Q_out814), // LUT general output
		.I0(Q_out813) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst815(
		.O(Q_out815), // LUT general output
		.I0(Q_out814) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst816(
		.O(Q_out816), // LUT general output
		.I0(Q_out815) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst817(
		.O(Q_out817), // LUT general output
		.I0(Q_out816) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst818(
		.O(Q_out818), // LUT general output
		.I0(Q_out817) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst819(
		.O(Q_out819), // LUT general output
		.I0(Q_out818) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst820(
		.O(Q_out820), // LUT general output
		.I0(Q_out819) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst821(
		.O(Q_out821), // LUT general output
		.I0(Q_out820) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst822(
		.O(Q_out822), // LUT general output
		.I0(Q_out821) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst823(
		.O(Q_out823), // LUT general output
		.I0(Q_out822) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst824(
		.O(Q_out824), // LUT general output
		.I0(Q_out823) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst825(
		.O(Q_out825), // LUT general output
		.I0(Q_out824) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst826(
		.O(Q_out826), // LUT general output
		.I0(Q_out825) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst827(
		.O(Q_out827), // LUT general output
		.I0(Q_out826) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst828(
		.O(Q_out828), // LUT general output
		.I0(Q_out827) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst829(
		.O(Q_out829), // LUT general output
		.I0(Q_out828) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst830(
		.O(Q_out830), // LUT general output
		.I0(Q_out829) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst831(
		.O(Q_out831), // LUT general output
		.I0(Q_out830) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst832(
		.O(Q_out832), // LUT general output
		.I0(Q_out831) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst833(
		.O(Q_out833), // LUT general output
		.I0(Q_out832) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst834(
		.O(Q_out834), // LUT general output
		.I0(Q_out833) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst835(
		.O(Q_out835), // LUT general output
		.I0(Q_out834) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst836(
		.O(Q_out836), // LUT general output
		.I0(Q_out835) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst837(
		.O(Q_out837), // LUT general output
		.I0(Q_out836) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst838(
		.O(Q_out838), // LUT general output
		.I0(Q_out837) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst839(
		.O(Q_out839), // LUT general output
		.I0(Q_out838) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst840(
		.O(Q_out840), // LUT general output
		.I0(Q_out839) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst841(
		.O(Q_out841), // LUT general output
		.I0(Q_out840) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst842(
		.O(Q_out842), // LUT general output
		.I0(Q_out841) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst843(
		.O(Q_out843), // LUT general output
		.I0(Q_out842) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst844(
		.O(Q_out844), // LUT general output
		.I0(Q_out843) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst845(
		.O(Q_out845), // LUT general output
		.I0(Q_out844) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst846(
		.O(Q_out846), // LUT general output
		.I0(Q_out845) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst847(
		.O(Q_out847), // LUT general output
		.I0(Q_out846) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst848(
		.O(Q_out848), // LUT general output
		.I0(Q_out847) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst849(
		.O(Q_out849), // LUT general output
		.I0(Q_out848) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst850(
		.O(Q_out850), // LUT general output
		.I0(Q_out849) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst851(
		.O(Q_out851), // LUT general output
		.I0(Q_out850) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst852(
		.O(Q_out852), // LUT general output
		.I0(Q_out851) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst853(
		.O(Q_out853), // LUT general output
		.I0(Q_out852) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst854(
		.O(Q_out854), // LUT general output
		.I0(Q_out853) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst855(
		.O(Q_out855), // LUT general output
		.I0(Q_out854) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst856(
		.O(Q_out856), // LUT general output
		.I0(Q_out855) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst857(
		.O(Q_out857), // LUT general output
		.I0(Q_out856) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst858(
		.O(Q_out858), // LUT general output
		.I0(Q_out857) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst859(
		.O(Q_out859), // LUT general output
		.I0(Q_out858) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst860(
		.O(Q_out860), // LUT general output
		.I0(Q_out859) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst861(
		.O(Q_out861), // LUT general output
		.I0(Q_out860) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst862(
		.O(Q_out862), // LUT general output
		.I0(Q_out861) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst863(
		.O(Q_out863), // LUT general output
		.I0(Q_out862) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst864(
		.O(Q_out864), // LUT general output
		.I0(Q_out863) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst865(
		.O(Q_out865), // LUT general output
		.I0(Q_out864) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst866(
		.O(Q_out866), // LUT general output
		.I0(Q_out865) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst867(
		.O(Q_out867), // LUT general output
		.I0(Q_out866) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst868(
		.O(Q_out868), // LUT general output
		.I0(Q_out867) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst869(
		.O(Q_out869), // LUT general output
		.I0(Q_out868) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst870(
		.O(Q_out870), // LUT general output
		.I0(Q_out869) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst871(
		.O(Q_out871), // LUT general output
		.I0(Q_out870) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst872(
		.O(Q_out872), // LUT general output
		.I0(Q_out871) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst873(
		.O(Q_out873), // LUT general output
		.I0(Q_out872) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst874(
		.O(Q_out874), // LUT general output
		.I0(Q_out873) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst875(
		.O(Q_out875), // LUT general output
		.I0(Q_out874) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst876(
		.O(Q_out876), // LUT general output
		.I0(Q_out875) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst877(
		.O(Q_out877), // LUT general output
		.I0(Q_out876) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst878(
		.O(Q_out878), // LUT general output
		.I0(Q_out877) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst879(
		.O(Q_out879), // LUT general output
		.I0(Q_out878) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst880(
		.O(Q_out880), // LUT general output
		.I0(Q_out879) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst881(
		.O(Q_out881), // LUT general output
		.I0(Q_out880) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst882(
		.O(Q_out882), // LUT general output
		.I0(Q_out881) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst883(
		.O(Q_out883), // LUT general output
		.I0(Q_out882) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst884(
		.O(Q_out884), // LUT general output
		.I0(Q_out883) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst885(
		.O(Q_out885), // LUT general output
		.I0(Q_out884) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst886(
		.O(Q_out886), // LUT general output
		.I0(Q_out885) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst887(
		.O(Q_out887), // LUT general output
		.I0(Q_out886) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst888(
		.O(Q_out888), // LUT general output
		.I0(Q_out887) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst889(
		.O(Q_out889), // LUT general output
		.I0(Q_out888) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst890(
		.O(Q_out890), // LUT general output
		.I0(Q_out889) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst891(
		.O(Q_out891), // LUT general output
		.I0(Q_out890) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst892(
		.O(Q_out892), // LUT general output
		.I0(Q_out891) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst893(
		.O(Q_out893), // LUT general output
		.I0(Q_out892) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst894(
		.O(Q_out894), // LUT general output
		.I0(Q_out893) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst895(
		.O(Q_out895), // LUT general output
		.I0(Q_out894) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst896(
		.O(Q_out896), // LUT general output
		.I0(Q_out895) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst897(
		.O(Q_out897), // LUT general output
		.I0(Q_out896) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst898(
		.O(Q_out898), // LUT general output
		.I0(Q_out897) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst899(
		.O(Q_out899), // LUT general output
		.I0(Q_out898) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst900(
		.O(Q_out900), // LUT general output
		.I0(Q_out899) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst901(
		.O(Q_out901), // LUT general output
		.I0(Q_out900) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst902(
		.O(Q_out902), // LUT general output
		.I0(Q_out901) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst903(
		.O(Q_out903), // LUT general output
		.I0(Q_out902) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst904(
		.O(Q_out904), // LUT general output
		.I0(Q_out903) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst905(
		.O(Q_out905), // LUT general output
		.I0(Q_out904) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst906(
		.O(Q_out906), // LUT general output
		.I0(Q_out905) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst907(
		.O(Q_out907), // LUT general output
		.I0(Q_out906) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst908(
		.O(Q_out908), // LUT general output
		.I0(Q_out907) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst909(
		.O(Q_out909), // LUT general output
		.I0(Q_out908) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst910(
		.O(Q_out910), // LUT general output
		.I0(Q_out909) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst911(
		.O(Q_out911), // LUT general output
		.I0(Q_out910) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst912(
		.O(Q_out912), // LUT general output
		.I0(Q_out911) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst913(
		.O(Q_out913), // LUT general output
		.I0(Q_out912) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst914(
		.O(Q_out914), // LUT general output
		.I0(Q_out913) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst915(
		.O(Q_out915), // LUT general output
		.I0(Q_out914) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst916(
		.O(Q_out916), // LUT general output
		.I0(Q_out915) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst917(
		.O(Q_out917), // LUT general output
		.I0(Q_out916) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst918(
		.O(Q_out918), // LUT general output
		.I0(Q_out917) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst919(
		.O(Q_out919), // LUT general output
		.I0(Q_out918) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst920(
		.O(Q_out920), // LUT general output
		.I0(Q_out919) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst921(
		.O(Q_out921), // LUT general output
		.I0(Q_out920) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst922(
		.O(Q_out922), // LUT general output
		.I0(Q_out921) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst923(
		.O(Q_out923), // LUT general output
		.I0(Q_out922) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst924(
		.O(Q_out924), // LUT general output
		.I0(Q_out923) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst925(
		.O(Q_out925), // LUT general output
		.I0(Q_out924) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst926(
		.O(Q_out926), // LUT general output
		.I0(Q_out925) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst927(
		.O(Q_out927), // LUT general output
		.I0(Q_out926) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst928(
		.O(Q_out928), // LUT general output
		.I0(Q_out927) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst929(
		.O(Q_out929), // LUT general output
		.I0(Q_out928) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst930(
		.O(Q_out930), // LUT general output
		.I0(Q_out929) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst931(
		.O(Q_out931), // LUT general output
		.I0(Q_out930) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst932(
		.O(Q_out932), // LUT general output
		.I0(Q_out931) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst933(
		.O(Q_out933), // LUT general output
		.I0(Q_out932) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst934(
		.O(Q_out934), // LUT general output
		.I0(Q_out933) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst935(
		.O(Q_out935), // LUT general output
		.I0(Q_out934) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst936(
		.O(Q_out936), // LUT general output
		.I0(Q_out935) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst937(
		.O(Q_out937), // LUT general output
		.I0(Q_out936) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst938(
		.O(Q_out938), // LUT general output
		.I0(Q_out937) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst939(
		.O(Q_out939), // LUT general output
		.I0(Q_out938) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst940(
		.O(Q_out940), // LUT general output
		.I0(Q_out939) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst941(
		.O(Q_out941), // LUT general output
		.I0(Q_out940) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst942(
		.O(Q_out942), // LUT general output
		.I0(Q_out941) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst943(
		.O(Q_out943), // LUT general output
		.I0(Q_out942) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst944(
		.O(Q_out944), // LUT general output
		.I0(Q_out943) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst945(
		.O(Q_out945), // LUT general output
		.I0(Q_out944) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst946(
		.O(Q_out946), // LUT general output
		.I0(Q_out945) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst947(
		.O(Q_out947), // LUT general output
		.I0(Q_out946) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst948(
		.O(Q_out948), // LUT general output
		.I0(Q_out947) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst949(
		.O(Q_out949), // LUT general output
		.I0(Q_out948) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst950(
		.O(Q_out950), // LUT general output
		.I0(Q_out949) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst951(
		.O(Q_out951), // LUT general output
		.I0(Q_out950) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst952(
		.O(Q_out952), // LUT general output
		.I0(Q_out951) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst953(
		.O(Q_out953), // LUT general output
		.I0(Q_out952) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst954(
		.O(Q_out954), // LUT general output
		.I0(Q_out953) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst955(
		.O(Q_out955), // LUT general output
		.I0(Q_out954) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst956(
		.O(Q_out956), // LUT general output
		.I0(Q_out955) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst957(
		.O(Q_out957), // LUT general output
		.I0(Q_out956) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst958(
		.O(Q_out958), // LUT general output
		.I0(Q_out957) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst959(
		.O(Q_out959), // LUT general output
		.I0(Q_out958) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst960(
		.O(Q_out960), // LUT general output
		.I0(Q_out959) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst961(
		.O(Q_out961), // LUT general output
		.I0(Q_out960) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst962(
		.O(Q_out962), // LUT general output
		.I0(Q_out961) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst963(
		.O(Q_out963), // LUT general output
		.I0(Q_out962) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst964(
		.O(Q_out964), // LUT general output
		.I0(Q_out963) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst965(
		.O(Q_out965), // LUT general output
		.I0(Q_out964) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst966(
		.O(Q_out966), // LUT general output
		.I0(Q_out965) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst967(
		.O(Q_out967), // LUT general output
		.I0(Q_out966) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst968(
		.O(Q_out968), // LUT general output
		.I0(Q_out967) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst969(
		.O(Q_out969), // LUT general output
		.I0(Q_out968) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst970(
		.O(Q_out970), // LUT general output
		.I0(Q_out969) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst971(
		.O(Q_out971), // LUT general output
		.I0(Q_out970) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst972(
		.O(Q_out972), // LUT general output
		.I0(Q_out971) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst973(
		.O(Q_out973), // LUT general output
		.I0(Q_out972) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst974(
		.O(Q_out974), // LUT general output
		.I0(Q_out973) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst975(
		.O(Q_out975), // LUT general output
		.I0(Q_out974) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst976(
		.O(Q_out976), // LUT general output
		.I0(Q_out975) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst977(
		.O(Q_out977), // LUT general output
		.I0(Q_out976) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst978(
		.O(Q_out978), // LUT general output
		.I0(Q_out977) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst979(
		.O(Q_out979), // LUT general output
		.I0(Q_out978) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst980(
		.O(Q_out980), // LUT general output
		.I0(Q_out979) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst981(
		.O(Q_out981), // LUT general output
		.I0(Q_out980) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst982(
		.O(Q_out982), // LUT general output
		.I0(Q_out981) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst983(
		.O(Q_out983), // LUT general output
		.I0(Q_out982) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst984(
		.O(Q_out984), // LUT general output
		.I0(Q_out983) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst985(
		.O(Q_out985), // LUT general output
		.I0(Q_out984) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst986(
		.O(Q_out986), // LUT general output
		.I0(Q_out985) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst987(
		.O(Q_out987), // LUT general output
		.I0(Q_out986) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst988(
		.O(Q_out988), // LUT general output
		.I0(Q_out987) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst989(
		.O(Q_out989), // LUT general output
		.I0(Q_out988) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst990(
		.O(Q_out990), // LUT general output
		.I0(Q_out989) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst991(
		.O(Q_out991), // LUT general output
		.I0(Q_out990) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst992(
		.O(Q_out992), // LUT general output
		.I0(Q_out991) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst993(
		.O(Q_out993), // LUT general output
		.I0(Q_out992) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst994(
		.O(Q_out994), // LUT general output
		.I0(Q_out993) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst995(
		.O(Q_out995), // LUT general output
		.I0(Q_out994) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst996(
		.O(Q_out996), // LUT general output
		.I0(Q_out995) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst997(
		.O(Q_out997), // LUT general output
		.I0(Q_out996) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst998(
		.O(Q_out998), // LUT general output
		.I0(Q_out997) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst999(
		.O(Q_out999), // LUT general output
		.I0(Q_out998) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1000(
		.O(Q_out1000), // LUT general output
		.I0(Q_out999) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1001(
		.O(Q_out1001), // LUT general output
		.I0(Q_out1000) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1002(
		.O(Q_out1002), // LUT general output
		.I0(Q_out1001) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1003(
		.O(Q_out1003), // LUT general output
		.I0(Q_out1002) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1004(
		.O(Q_out1004), // LUT general output
		.I0(Q_out1003) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1005(
		.O(Q_out1005), // LUT general output
		.I0(Q_out1004) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1006(
		.O(Q_out1006), // LUT general output
		.I0(Q_out1005) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1007(
		.O(Q_out1007), // LUT general output
		.I0(Q_out1006) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1008(
		.O(Q_out1008), // LUT general output
		.I0(Q_out1007) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1009(
		.O(Q_out1009), // LUT general output
		.I0(Q_out1008) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1010(
		.O(Q_out1010), // LUT general output
		.I0(Q_out1009) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1011(
		.O(Q_out1011), // LUT general output
		.I0(Q_out1010) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1012(
		.O(Q_out1012), // LUT general output
		.I0(Q_out1011) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1013(
		.O(Q_out1013), // LUT general output
		.I0(Q_out1012) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1014(
		.O(Q_out1014), // LUT general output
		.I0(Q_out1013) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1015(
		.O(Q_out1015), // LUT general output
		.I0(Q_out1014) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1016(
		.O(Q_out1016), // LUT general output
		.I0(Q_out1015) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1017(
		.O(Q_out1017), // LUT general output
		.I0(Q_out1016) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1018(
		.O(Q_out1018), // LUT general output
		.I0(Q_out1017) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1019(
		.O(Q_out1019), // LUT general output
		.I0(Q_out1018) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1020(
		.O(Q_out1020), // LUT general output
		.I0(Q_out1019) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1021(
		.O(Q_out1021), // LUT general output
		.I0(Q_out1020) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1022(
		.O(Q_out1022), // LUT general output
		.I0(Q_out1021) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1023(
		.O(Q_out1023), // LUT general output
		.I0(Q_out1022) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1024(
		.O(Q_out1024), // LUT general output
		.I0(Q_out1023) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1025(
		.O(Q_out1025), // LUT general output
		.I0(Q_out1024) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1026(
		.O(Q_out1026), // LUT general output
		.I0(Q_out1025) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1027(
		.O(Q_out1027), // LUT general output
		.I0(Q_out1026) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1028(
		.O(Q_out1028), // LUT general output
		.I0(Q_out1027) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1029(
		.O(Q_out1029), // LUT general output
		.I0(Q_out1028) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1030(
		.O(Q_out1030), // LUT general output
		.I0(Q_out1029) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1031(
		.O(Q_out1031), // LUT general output
		.I0(Q_out1030) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1032(
		.O(Q_out1032), // LUT general output
		.I0(Q_out1031) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1033(
		.O(Q_out1033), // LUT general output
		.I0(Q_out1032) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1034(
		.O(Q_out1034), // LUT general output
		.I0(Q_out1033) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1035(
		.O(Q_out1035), // LUT general output
		.I0(Q_out1034) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1036(
		.O(Q_out1036), // LUT general output
		.I0(Q_out1035) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1037(
		.O(Q_out1037), // LUT general output
		.I0(Q_out1036) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1038(
		.O(Q_out1038), // LUT general output
		.I0(Q_out1037) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1039(
		.O(Q_out1039), // LUT general output
		.I0(Q_out1038) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1040(
		.O(Q_out1040), // LUT general output
		.I0(Q_out1039) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1041(
		.O(Q_out1041), // LUT general output
		.I0(Q_out1040) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1042(
		.O(Q_out1042), // LUT general output
		.I0(Q_out1041) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1043(
		.O(Q_out1043), // LUT general output
		.I0(Q_out1042) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1044(
		.O(Q_out1044), // LUT general output
		.I0(Q_out1043) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1045(
		.O(Q_out1045), // LUT general output
		.I0(Q_out1044) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1046(
		.O(Q_out1046), // LUT general output
		.I0(Q_out1045) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1047(
		.O(Q_out1047), // LUT general output
		.I0(Q_out1046) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1048(
		.O(Q_out1048), // LUT general output
		.I0(Q_out1047) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1049(
		.O(Q_out1049), // LUT general output
		.I0(Q_out1048) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1050(
		.O(Q_out1050), // LUT general output
		.I0(Q_out1049) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1051(
		.O(Q_out1051), // LUT general output
		.I0(Q_out1050) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1052(
		.O(Q_out1052), // LUT general output
		.I0(Q_out1051) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1053(
		.O(Q_out1053), // LUT general output
		.I0(Q_out1052) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1054(
		.O(Q_out1054), // LUT general output
		.I0(Q_out1053) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1055(
		.O(Q_out1055), // LUT general output
		.I0(Q_out1054) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1056(
		.O(Q_out1056), // LUT general output
		.I0(Q_out1055) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1057(
		.O(Q_out1057), // LUT general output
		.I0(Q_out1056) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1058(
		.O(Q_out1058), // LUT general output
		.I0(Q_out1057) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1059(
		.O(Q_out1059), // LUT general output
		.I0(Q_out1058) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1060(
		.O(Q_out1060), // LUT general output
		.I0(Q_out1059) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1061(
		.O(Q_out1061), // LUT general output
		.I0(Q_out1060) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1062(
		.O(Q_out1062), // LUT general output
		.I0(Q_out1061) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1063(
		.O(Q_out1063), // LUT general output
		.I0(Q_out1062) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1064(
		.O(Q_out1064), // LUT general output
		.I0(Q_out1063) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1065(
		.O(Q_out1065), // LUT general output
		.I0(Q_out1064) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1066(
		.O(Q_out1066), // LUT general output
		.I0(Q_out1065) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1067(
		.O(Q_out1067), // LUT general output
		.I0(Q_out1066) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1068(
		.O(Q_out1068), // LUT general output
		.I0(Q_out1067) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1069(
		.O(Q_out1069), // LUT general output
		.I0(Q_out1068) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1070(
		.O(Q_out1070), // LUT general output
		.I0(Q_out1069) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1071(
		.O(Q_out1071), // LUT general output
		.I0(Q_out1070) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1072(
		.O(Q_out1072), // LUT general output
		.I0(Q_out1071) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1073(
		.O(Q_out1073), // LUT general output
		.I0(Q_out1072) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1074(
		.O(Q_out1074), // LUT general output
		.I0(Q_out1073) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1075(
		.O(Q_out1075), // LUT general output
		.I0(Q_out1074) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1076(
		.O(Q_out1076), // LUT general output
		.I0(Q_out1075) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1077(
		.O(Q_out1077), // LUT general output
		.I0(Q_out1076) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1078(
		.O(Q_out1078), // LUT general output
		.I0(Q_out1077) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1079(
		.O(Q_out1079), // LUT general output
		.I0(Q_out1078) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1080(
		.O(Q_out1080), // LUT general output
		.I0(Q_out1079) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1081(
		.O(Q_out1081), // LUT general output
		.I0(Q_out1080) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1082(
		.O(Q_out1082), // LUT general output
		.I0(Q_out1081) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1083(
		.O(Q_out1083), // LUT general output
		.I0(Q_out1082) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1084(
		.O(Q_out1084), // LUT general output
		.I0(Q_out1083) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1085(
		.O(Q_out1085), // LUT general output
		.I0(Q_out1084) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1086(
		.O(Q_out1086), // LUT general output
		.I0(Q_out1085) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1087(
		.O(Q_out1087), // LUT general output
		.I0(Q_out1086) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1088(
		.O(Q_out1088), // LUT general output
		.I0(Q_out1087) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1089(
		.O(Q_out1089), // LUT general output
		.I0(Q_out1088) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1090(
		.O(Q_out1090), // LUT general output
		.I0(Q_out1089) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1091(
		.O(Q_out1091), // LUT general output
		.I0(Q_out1090) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1092(
		.O(Q_out1092), // LUT general output
		.I0(Q_out1091) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1093(
		.O(Q_out1093), // LUT general output
		.I0(Q_out1092) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1094(
		.O(Q_out1094), // LUT general output
		.I0(Q_out1093) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1095(
		.O(Q_out1095), // LUT general output
		.I0(Q_out1094) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1096(
		.O(Q_out1096), // LUT general output
		.I0(Q_out1095) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1097(
		.O(Q_out1097), // LUT general output
		.I0(Q_out1096) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1098(
		.O(Q_out1098), // LUT general output
		.I0(Q_out1097) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1099(
		.O(Q_out1099), // LUT general output
		.I0(Q_out1098) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1100(
		.O(Q_out1100), // LUT general output
		.I0(Q_out1099) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1101(
		.O(Q_out1101), // LUT general output
		.I0(Q_out1100) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1102(
		.O(Q_out1102), // LUT general output
		.I0(Q_out1101) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1103(
		.O(Q_out1103), // LUT general output
		.I0(Q_out1102) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1104(
		.O(Q_out1104), // LUT general output
		.I0(Q_out1103) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1105(
		.O(Q_out1105), // LUT general output
		.I0(Q_out1104) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1106(
		.O(Q_out1106), // LUT general output
		.I0(Q_out1105) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1107(
		.O(Q_out1107), // LUT general output
		.I0(Q_out1106) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1108(
		.O(Q_out1108), // LUT general output
		.I0(Q_out1107) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1109(
		.O(Q_out1109), // LUT general output
		.I0(Q_out1108) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1110(
		.O(Q_out1110), // LUT general output
		.I0(Q_out1109) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1111(
		.O(Q_out1111), // LUT general output
		.I0(Q_out1110) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1112(
		.O(Q_out1112), // LUT general output
		.I0(Q_out1111) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1113(
		.O(Q_out1113), // LUT general output
		.I0(Q_out1112) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1114(
		.O(Q_out1114), // LUT general output
		.I0(Q_out1113) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1115(
		.O(Q_out1115), // LUT general output
		.I0(Q_out1114) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1116(
		.O(Q_out1116), // LUT general output
		.I0(Q_out1115) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1117(
		.O(Q_out1117), // LUT general output
		.I0(Q_out1116) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1118(
		.O(Q_out1118), // LUT general output
		.I0(Q_out1117) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1119(
		.O(Q_out1119), // LUT general output
		.I0(Q_out1118) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1120(
		.O(Q_out1120), // LUT general output
		.I0(Q_out1119) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1121(
		.O(Q_out1121), // LUT general output
		.I0(Q_out1120) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1122(
		.O(Q_out1122), // LUT general output
		.I0(Q_out1121) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1123(
		.O(Q_out1123), // LUT general output
		.I0(Q_out1122) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1124(
		.O(Q_out1124), // LUT general output
		.I0(Q_out1123) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1125(
		.O(Q_out1125), // LUT general output
		.I0(Q_out1124) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1126(
		.O(Q_out1126), // LUT general output
		.I0(Q_out1125) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1127(
		.O(Q_out1127), // LUT general output
		.I0(Q_out1126) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1128(
		.O(Q_out1128), // LUT general output
		.I0(Q_out1127) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1129(
		.O(Q_out1129), // LUT general output
		.I0(Q_out1128) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1130(
		.O(Q_out1130), // LUT general output
		.I0(Q_out1129) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1131(
		.O(Q_out1131), // LUT general output
		.I0(Q_out1130) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1132(
		.O(Q_out1132), // LUT general output
		.I0(Q_out1131) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1133(
		.O(Q_out1133), // LUT general output
		.I0(Q_out1132) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1134(
		.O(Q_out1134), // LUT general output
		.I0(Q_out1133) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1135(
		.O(Q_out1135), // LUT general output
		.I0(Q_out1134) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1136(
		.O(Q_out1136), // LUT general output
		.I0(Q_out1135) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1137(
		.O(Q_out1137), // LUT general output
		.I0(Q_out1136) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1138(
		.O(Q_out1138), // LUT general output
		.I0(Q_out1137) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1139(
		.O(Q_out1139), // LUT general output
		.I0(Q_out1138) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1140(
		.O(Q_out1140), // LUT general output
		.I0(Q_out1139) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1141(
		.O(Q_out1141), // LUT general output
		.I0(Q_out1140) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1142(
		.O(Q_out1142), // LUT general output
		.I0(Q_out1141) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1143(
		.O(Q_out1143), // LUT general output
		.I0(Q_out1142) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1144(
		.O(Q_out1144), // LUT general output
		.I0(Q_out1143) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1145(
		.O(Q_out1145), // LUT general output
		.I0(Q_out1144) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1146(
		.O(Q_out1146), // LUT general output
		.I0(Q_out1145) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1147(
		.O(Q_out1147), // LUT general output
		.I0(Q_out1146) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1148(
		.O(Q_out1148), // LUT general output
		.I0(Q_out1147) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1149(
		.O(Q_out1149), // LUT general output
		.I0(Q_out1148) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1150(
		.O(Q_out1150), // LUT general output
		.I0(Q_out1149) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1151(
		.O(Q_out1151), // LUT general output
		.I0(Q_out1150) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1152(
		.O(Q_out1152), // LUT general output
		.I0(Q_out1151) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1153(
		.O(Q_out1153), // LUT general output
		.I0(Q_out1152) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1154(
		.O(Q_out1154), // LUT general output
		.I0(Q_out1153) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1155(
		.O(Q_out1155), // LUT general output
		.I0(Q_out1154) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1156(
		.O(Q_out1156), // LUT general output
		.I0(Q_out1155) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1157(
		.O(Q_out1157), // LUT general output
		.I0(Q_out1156) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1158(
		.O(Q_out1158), // LUT general output
		.I0(Q_out1157) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1159(
		.O(Q_out1159), // LUT general output
		.I0(Q_out1158) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1160(
		.O(Q_out1160), // LUT general output
		.I0(Q_out1159) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1161(
		.O(Q_out1161), // LUT general output
		.I0(Q_out1160) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1162(
		.O(Q_out1162), // LUT general output
		.I0(Q_out1161) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1163(
		.O(Q_out1163), // LUT general output
		.I0(Q_out1162) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1164(
		.O(Q_out1164), // LUT general output
		.I0(Q_out1163) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1165(
		.O(Q_out1165), // LUT general output
		.I0(Q_out1164) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1166(
		.O(Q_out1166), // LUT general output
		.I0(Q_out1165) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1167(
		.O(Q_out1167), // LUT general output
		.I0(Q_out1166) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1168(
		.O(Q_out1168), // LUT general output
		.I0(Q_out1167) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1169(
		.O(Q_out1169), // LUT general output
		.I0(Q_out1168) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1170(
		.O(Q_out1170), // LUT general output
		.I0(Q_out1169) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1171(
		.O(Q_out1171), // LUT general output
		.I0(Q_out1170) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1172(
		.O(Q_out1172), // LUT general output
		.I0(Q_out1171) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1173(
		.O(Q_out1173), // LUT general output
		.I0(Q_out1172) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1174(
		.O(Q_out1174), // LUT general output
		.I0(Q_out1173) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1175(
		.O(Q_out1175), // LUT general output
		.I0(Q_out1174) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1176(
		.O(Q_out1176), // LUT general output
		.I0(Q_out1175) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1177(
		.O(Q_out1177), // LUT general output
		.I0(Q_out1176) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1178(
		.O(Q_out1178), // LUT general output
		.I0(Q_out1177) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1179(
		.O(Q_out1179), // LUT general output
		.I0(Q_out1178) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1180(
		.O(Q_out1180), // LUT general output
		.I0(Q_out1179) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1181(
		.O(Q_out1181), // LUT general output
		.I0(Q_out1180) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1182(
		.O(Q_out1182), // LUT general output
		.I0(Q_out1181) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1183(
		.O(Q_out1183), // LUT general output
		.I0(Q_out1182) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1184(
		.O(Q_out1184), // LUT general output
		.I0(Q_out1183) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1185(
		.O(Q_out1185), // LUT general output
		.I0(Q_out1184) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1186(
		.O(Q_out1186), // LUT general output
		.I0(Q_out1185) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1187(
		.O(Q_out1187), // LUT general output
		.I0(Q_out1186) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1188(
		.O(Q_out1188), // LUT general output
		.I0(Q_out1187) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1189(
		.O(Q_out1189), // LUT general output
		.I0(Q_out1188) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1190(
		.O(Q_out1190), // LUT general output
		.I0(Q_out1189) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1191(
		.O(Q_out1191), // LUT general output
		.I0(Q_out1190) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1192(
		.O(Q_out1192), // LUT general output
		.I0(Q_out1191) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1193(
		.O(Q_out1193), // LUT general output
		.I0(Q_out1192) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1194(
		.O(Q_out1194), // LUT general output
		.I0(Q_out1193) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1195(
		.O(Q_out1195), // LUT general output
		.I0(Q_out1194) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1196(
		.O(Q_out1196), // LUT general output
		.I0(Q_out1195) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1197(
		.O(Q_out1197), // LUT general output
		.I0(Q_out1196) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1198(
		.O(Q_out1198), // LUT general output
		.I0(Q_out1197) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1199(
		.O(Q_out1199), // LUT general output
		.I0(Q_out1198) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1200(
		.O(Q_out1200), // LUT general output
		.I0(Q_out1199) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1201(
		.O(Q_out1201), // LUT general output
		.I0(Q_out1200) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1202(
		.O(Q_out1202), // LUT general output
		.I0(Q_out1201) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1203(
		.O(Q_out1203), // LUT general output
		.I0(Q_out1202) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1204(
		.O(Q_out1204), // LUT general output
		.I0(Q_out1203) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1205(
		.O(Q_out1205), // LUT general output
		.I0(Q_out1204) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1206(
		.O(Q_out1206), // LUT general output
		.I0(Q_out1205) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1207(
		.O(Q_out1207), // LUT general output
		.I0(Q_out1206) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1208(
		.O(Q_out1208), // LUT general output
		.I0(Q_out1207) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1209(
		.O(Q_out1209), // LUT general output
		.I0(Q_out1208) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1210(
		.O(Q_out1210), // LUT general output
		.I0(Q_out1209) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1211(
		.O(Q_out1211), // LUT general output
		.I0(Q_out1210) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1212(
		.O(Q_out1212), // LUT general output
		.I0(Q_out1211) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1213(
		.O(Q_out1213), // LUT general output
		.I0(Q_out1212) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1214(
		.O(Q_out1214), // LUT general output
		.I0(Q_out1213) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1215(
		.O(Q_out1215), // LUT general output
		.I0(Q_out1214) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1216(
		.O(Q_out1216), // LUT general output
		.I0(Q_out1215) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1217(
		.O(Q_out1217), // LUT general output
		.I0(Q_out1216) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1218(
		.O(Q_out1218), // LUT general output
		.I0(Q_out1217) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1219(
		.O(Q_out1219), // LUT general output
		.I0(Q_out1218) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1220(
		.O(Q_out1220), // LUT general output
		.I0(Q_out1219) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1221(
		.O(Q_out1221), // LUT general output
		.I0(Q_out1220) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1222(
		.O(Q_out1222), // LUT general output
		.I0(Q_out1221) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1223(
		.O(Q_out1223), // LUT general output
		.I0(Q_out1222) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1224(
		.O(Q_out1224), // LUT general output
		.I0(Q_out1223) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1225(
		.O(Q_out1225), // LUT general output
		.I0(Q_out1224) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1226(
		.O(Q_out1226), // LUT general output
		.I0(Q_out1225) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1227(
		.O(Q_out1227), // LUT general output
		.I0(Q_out1226) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1228(
		.O(Q_out1228), // LUT general output
		.I0(Q_out1227) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1229(
		.O(Q_out1229), // LUT general output
		.I0(Q_out1228) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1230(
		.O(Q_out1230), // LUT general output
		.I0(Q_out1229) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1231(
		.O(Q_out1231), // LUT general output
		.I0(Q_out1230) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1232(
		.O(Q_out1232), // LUT general output
		.I0(Q_out1231) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1233(
		.O(Q_out1233), // LUT general output
		.I0(Q_out1232) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1234(
		.O(Q_out1234), // LUT general output
		.I0(Q_out1233) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1235(
		.O(Q_out1235), // LUT general output
		.I0(Q_out1234) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1236(
		.O(Q_out1236), // LUT general output
		.I0(Q_out1235) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1237(
		.O(Q_out1237), // LUT general output
		.I0(Q_out1236) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1238(
		.O(Q_out1238), // LUT general output
		.I0(Q_out1237) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1239(
		.O(Q_out1239), // LUT general output
		.I0(Q_out1238) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1240(
		.O(Q_out1240), // LUT general output
		.I0(Q_out1239) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1241(
		.O(Q_out1241), // LUT general output
		.I0(Q_out1240) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1242(
		.O(Q_out1242), // LUT general output
		.I0(Q_out1241) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1243(
		.O(Q_out1243), // LUT general output
		.I0(Q_out1242) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1244(
		.O(Q_out1244), // LUT general output
		.I0(Q_out1243) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1245(
		.O(Q_out1245), // LUT general output
		.I0(Q_out1244) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1246(
		.O(Q_out1246), // LUT general output
		.I0(Q_out1245) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1247(
		.O(Q_out1247), // LUT general output
		.I0(Q_out1246) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1248(
		.O(Q_out1248), // LUT general output
		.I0(Q_out1247) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1249(
		.O(Q_out1249), // LUT general output
		.I0(Q_out1248) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1250(
		.O(Q_out1250), // LUT general output
		.I0(Q_out1249) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1251(
		.O(Q_out1251), // LUT general output
		.I0(Q_out1250) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1252(
		.O(Q_out1252), // LUT general output
		.I0(Q_out1251) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1253(
		.O(Q_out1253), // LUT general output
		.I0(Q_out1252) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1254(
		.O(Q_out1254), // LUT general output
		.I0(Q_out1253) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1255(
		.O(Q_out1255), // LUT general output
		.I0(Q_out1254) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1256(
		.O(Q_out1256), // LUT general output
		.I0(Q_out1255) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1257(
		.O(Q_out1257), // LUT general output
		.I0(Q_out1256) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1258(
		.O(Q_out1258), // LUT general output
		.I0(Q_out1257) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1259(
		.O(Q_out1259), // LUT general output
		.I0(Q_out1258) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1260(
		.O(Q_out1260), // LUT general output
		.I0(Q_out1259) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1261(
		.O(Q_out1261), // LUT general output
		.I0(Q_out1260) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1262(
		.O(Q_out1262), // LUT general output
		.I0(Q_out1261) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1263(
		.O(Q_out1263), // LUT general output
		.I0(Q_out1262) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1264(
		.O(Q_out1264), // LUT general output
		.I0(Q_out1263) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1265(
		.O(Q_out1265), // LUT general output
		.I0(Q_out1264) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1266(
		.O(Q_out1266), // LUT general output
		.I0(Q_out1265) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1267(
		.O(Q_out1267), // LUT general output
		.I0(Q_out1266) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1268(
		.O(Q_out1268), // LUT general output
		.I0(Q_out1267) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1269(
		.O(Q_out1269), // LUT general output
		.I0(Q_out1268) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1270(
		.O(Q_out1270), // LUT general output
		.I0(Q_out1269) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1271(
		.O(Q_out1271), // LUT general output
		.I0(Q_out1270) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1272(
		.O(Q_out1272), // LUT general output
		.I0(Q_out1271) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1273(
		.O(Q_out1273), // LUT general output
		.I0(Q_out1272) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1274(
		.O(Q_out1274), // LUT general output
		.I0(Q_out1273) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1275(
		.O(Q_out1275), // LUT general output
		.I0(Q_out1274) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1276(
		.O(Q_out1276), // LUT general output
		.I0(Q_out1275) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1277(
		.O(Q_out1277), // LUT general output
		.I0(Q_out1276) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1278(
		.O(Q_out1278), // LUT general output
		.I0(Q_out1277) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1279(
		.O(Q_out1279), // LUT general output
		.I0(Q_out1278) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1280(
		.O(Q_out1280), // LUT general output
		.I0(Q_out1279) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1281(
		.O(Q_out1281), // LUT general output
		.I0(Q_out1280) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1282(
		.O(Q_out1282), // LUT general output
		.I0(Q_out1281) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1283(
		.O(Q_out1283), // LUT general output
		.I0(Q_out1282) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1284(
		.O(Q_out1284), // LUT general output
		.I0(Q_out1283) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1285(
		.O(Q_out1285), // LUT general output
		.I0(Q_out1284) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1286(
		.O(Q_out1286), // LUT general output
		.I0(Q_out1285) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1287(
		.O(Q_out1287), // LUT general output
		.I0(Q_out1286) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1288(
		.O(Q_out1288), // LUT general output
		.I0(Q_out1287) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1289(
		.O(Q_out1289), // LUT general output
		.I0(Q_out1288) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1290(
		.O(Q_out1290), // LUT general output
		.I0(Q_out1289) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1291(
		.O(Q_out1291), // LUT general output
		.I0(Q_out1290) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1292(
		.O(Q_out1292), // LUT general output
		.I0(Q_out1291) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1293(
		.O(Q_out1293), // LUT general output
		.I0(Q_out1292) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1294(
		.O(Q_out1294), // LUT general output
		.I0(Q_out1293) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1295(
		.O(Q_out1295), // LUT general output
		.I0(Q_out1294) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1296(
		.O(Q_out1296), // LUT general output
		.I0(Q_out1295) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1297(
		.O(Q_out1297), // LUT general output
		.I0(Q_out1296) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1298(
		.O(Q_out1298), // LUT general output
		.I0(Q_out1297) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1299(
		.O(Q_out1299), // LUT general output
		.I0(Q_out1298) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1300(
		.O(Q_out1300), // LUT general output
		.I0(Q_out1299) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1301(
		.O(Q_out1301), // LUT general output
		.I0(Q_out1300) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1302(
		.O(Q_out1302), // LUT general output
		.I0(Q_out1301) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1303(
		.O(Q_out1303), // LUT general output
		.I0(Q_out1302) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1304(
		.O(Q_out1304), // LUT general output
		.I0(Q_out1303) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1305(
		.O(Q_out1305), // LUT general output
		.I0(Q_out1304) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1306(
		.O(Q_out1306), // LUT general output
		.I0(Q_out1305) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1307(
		.O(Q_out1307), // LUT general output
		.I0(Q_out1306) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1308(
		.O(Q_out1308), // LUT general output
		.I0(Q_out1307) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1309(
		.O(Q_out1309), // LUT general output
		.I0(Q_out1308) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1310(
		.O(Q_out1310), // LUT general output
		.I0(Q_out1309) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1311(
		.O(Q_out1311), // LUT general output
		.I0(Q_out1310) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1312(
		.O(Q_out1312), // LUT general output
		.I0(Q_out1311) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1313(
		.O(Q_out1313), // LUT general output
		.I0(Q_out1312) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1314(
		.O(Q_out1314), // LUT general output
		.I0(Q_out1313) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1315(
		.O(Q_out1315), // LUT general output
		.I0(Q_out1314) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1316(
		.O(Q_out1316), // LUT general output
		.I0(Q_out1315) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1317(
		.O(Q_out1317), // LUT general output
		.I0(Q_out1316) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1318(
		.O(Q_out1318), // LUT general output
		.I0(Q_out1317) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1319(
		.O(Q_out1319), // LUT general output
		.I0(Q_out1318) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1320(
		.O(Q_out1320), // LUT general output
		.I0(Q_out1319) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1321(
		.O(Q_out1321), // LUT general output
		.I0(Q_out1320) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1322(
		.O(Q_out1322), // LUT general output
		.I0(Q_out1321) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1323(
		.O(Q_out1323), // LUT general output
		.I0(Q_out1322) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1324(
		.O(Q_out1324), // LUT general output
		.I0(Q_out1323) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1325(
		.O(Q_out1325), // LUT general output
		.I0(Q_out1324) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1326(
		.O(Q_out1326), // LUT general output
		.I0(Q_out1325) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1327(
		.O(Q_out1327), // LUT general output
		.I0(Q_out1326) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1328(
		.O(Q_out1328), // LUT general output
		.I0(Q_out1327) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1329(
		.O(Q_out1329), // LUT general output
		.I0(Q_out1328) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1330(
		.O(Q_out1330), // LUT general output
		.I0(Q_out1329) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1331(
		.O(Q_out1331), // LUT general output
		.I0(Q_out1330) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1332(
		.O(Q_out1332), // LUT general output
		.I0(Q_out1331) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1333(
		.O(Q_out1333), // LUT general output
		.I0(Q_out1332) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1334(
		.O(Q_out1334), // LUT general output
		.I0(Q_out1333) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1335(
		.O(Q_out1335), // LUT general output
		.I0(Q_out1334) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1336(
		.O(Q_out1336), // LUT general output
		.I0(Q_out1335) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1337(
		.O(Q_out1337), // LUT general output
		.I0(Q_out1336) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1338(
		.O(Q_out1338), // LUT general output
		.I0(Q_out1337) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1339(
		.O(Q_out1339), // LUT general output
		.I0(Q_out1338) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1340(
		.O(Q_out1340), // LUT general output
		.I0(Q_out1339) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1341(
		.O(Q_out1341), // LUT general output
		.I0(Q_out1340) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1342(
		.O(Q_out1342), // LUT general output
		.I0(Q_out1341) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1343(
		.O(Q_out1343), // LUT general output
		.I0(Q_out1342) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1344(
		.O(Q_out1344), // LUT general output
		.I0(Q_out1343) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1345(
		.O(Q_out1345), // LUT general output
		.I0(Q_out1344) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1346(
		.O(Q_out1346), // LUT general output
		.I0(Q_out1345) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1347(
		.O(Q_out1347), // LUT general output
		.I0(Q_out1346) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1348(
		.O(Q_out1348), // LUT general output
		.I0(Q_out1347) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1349(
		.O(Q_out1349), // LUT general output
		.I0(Q_out1348) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1350(
		.O(Q_out1350), // LUT general output
		.I0(Q_out1349) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1351(
		.O(Q_out1351), // LUT general output
		.I0(Q_out1350) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1352(
		.O(Q_out1352), // LUT general output
		.I0(Q_out1351) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1353(
		.O(Q_out1353), // LUT general output
		.I0(Q_out1352) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1354(
		.O(Q_out1354), // LUT general output
		.I0(Q_out1353) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1355(
		.O(Q_out1355), // LUT general output
		.I0(Q_out1354) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1356(
		.O(Q_out1356), // LUT general output
		.I0(Q_out1355) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1357(
		.O(Q_out1357), // LUT general output
		.I0(Q_out1356) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1358(
		.O(Q_out1358), // LUT general output
		.I0(Q_out1357) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1359(
		.O(Q_out1359), // LUT general output
		.I0(Q_out1358) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1360(
		.O(Q_out1360), // LUT general output
		.I0(Q_out1359) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1361(
		.O(Q_out1361), // LUT general output
		.I0(Q_out1360) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1362(
		.O(Q_out1362), // LUT general output
		.I0(Q_out1361) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1363(
		.O(Q_out1363), // LUT general output
		.I0(Q_out1362) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1364(
		.O(Q_out1364), // LUT general output
		.I0(Q_out1363) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1365(
		.O(Q_out1365), // LUT general output
		.I0(Q_out1364) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1366(
		.O(Q_out1366), // LUT general output
		.I0(Q_out1365) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1367(
		.O(Q_out1367), // LUT general output
		.I0(Q_out1366) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1368(
		.O(Q_out1368), // LUT general output
		.I0(Q_out1367) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1369(
		.O(Q_out1369), // LUT general output
		.I0(Q_out1368) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1370(
		.O(Q_out1370), // LUT general output
		.I0(Q_out1369) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1371(
		.O(Q_out1371), // LUT general output
		.I0(Q_out1370) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1372(
		.O(Q_out1372), // LUT general output
		.I0(Q_out1371) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1373(
		.O(Q_out1373), // LUT general output
		.I0(Q_out1372) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1374(
		.O(Q_out1374), // LUT general output
		.I0(Q_out1373) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1375(
		.O(Q_out1375), // LUT general output
		.I0(Q_out1374) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1376(
		.O(Q_out1376), // LUT general output
		.I0(Q_out1375) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1377(
		.O(Q_out1377), // LUT general output
		.I0(Q_out1376) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1378(
		.O(Q_out1378), // LUT general output
		.I0(Q_out1377) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1379(
		.O(Q_out1379), // LUT general output
		.I0(Q_out1378) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1380(
		.O(Q_out1380), // LUT general output
		.I0(Q_out1379) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1381(
		.O(Q_out1381), // LUT general output
		.I0(Q_out1380) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1382(
		.O(Q_out1382), // LUT general output
		.I0(Q_out1381) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1383(
		.O(Q_out1383), // LUT general output
		.I0(Q_out1382) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1384(
		.O(Q_out1384), // LUT general output
		.I0(Q_out1383) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1385(
		.O(Q_out1385), // LUT general output
		.I0(Q_out1384) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1386(
		.O(Q_out1386), // LUT general output
		.I0(Q_out1385) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1387(
		.O(Q_out1387), // LUT general output
		.I0(Q_out1386) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1388(
		.O(Q_out1388), // LUT general output
		.I0(Q_out1387) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1389(
		.O(Q_out1389), // LUT general output
		.I0(Q_out1388) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1390(
		.O(Q_out1390), // LUT general output
		.I0(Q_out1389) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1391(
		.O(Q_out1391), // LUT general output
		.I0(Q_out1390) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1392(
		.O(Q_out1392), // LUT general output
		.I0(Q_out1391) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1393(
		.O(Q_out1393), // LUT general output
		.I0(Q_out1392) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1394(
		.O(Q_out1394), // LUT general output
		.I0(Q_out1393) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1395(
		.O(Q_out1395), // LUT general output
		.I0(Q_out1394) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1396(
		.O(Q_out1396), // LUT general output
		.I0(Q_out1395) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1397(
		.O(Q_out1397), // LUT general output
		.I0(Q_out1396) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1398(
		.O(Q_out1398), // LUT general output
		.I0(Q_out1397) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1399(
		.O(Q_out1399), // LUT general output
		.I0(Q_out1398) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1400(
		.O(Q_out1400), // LUT general output
		.I0(Q_out1399) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1401(
		.O(Q_out1401), // LUT general output
		.I0(Q_out1400) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1402(
		.O(Q_out1402), // LUT general output
		.I0(Q_out1401) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1403(
		.O(Q_out1403), // LUT general output
		.I0(Q_out1402) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1404(
		.O(Q_out1404), // LUT general output
		.I0(Q_out1403) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1405(
		.O(Q_out1405), // LUT general output
		.I0(Q_out1404) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1406(
		.O(Q_out1406), // LUT general output
		.I0(Q_out1405) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1407(
		.O(Q_out1407), // LUT general output
		.I0(Q_out1406) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1408(
		.O(Q_out1408), // LUT general output
		.I0(Q_out1407) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1409(
		.O(Q_out1409), // LUT general output
		.I0(Q_out1408) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1410(
		.O(Q_out1410), // LUT general output
		.I0(Q_out1409) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1411(
		.O(Q_out1411), // LUT general output
		.I0(Q_out1410) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1412(
		.O(Q_out1412), // LUT general output
		.I0(Q_out1411) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1413(
		.O(Q_out1413), // LUT general output
		.I0(Q_out1412) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1414(
		.O(Q_out1414), // LUT general output
		.I0(Q_out1413) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1415(
		.O(Q_out1415), // LUT general output
		.I0(Q_out1414) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1416(
		.O(Q_out1416), // LUT general output
		.I0(Q_out1415) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1417(
		.O(Q_out1417), // LUT general output
		.I0(Q_out1416) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1418(
		.O(Q_out1418), // LUT general output
		.I0(Q_out1417) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1419(
		.O(Q_out1419), // LUT general output
		.I0(Q_out1418) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1420(
		.O(Q_out1420), // LUT general output
		.I0(Q_out1419) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1421(
		.O(Q_out1421), // LUT general output
		.I0(Q_out1420) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1422(
		.O(Q_out1422), // LUT general output
		.I0(Q_out1421) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1423(
		.O(Q_out1423), // LUT general output
		.I0(Q_out1422) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1424(
		.O(Q_out1424), // LUT general output
		.I0(Q_out1423) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1425(
		.O(Q_out1425), // LUT general output
		.I0(Q_out1424) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1426(
		.O(Q_out1426), // LUT general output
		.I0(Q_out1425) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1427(
		.O(Q_out1427), // LUT general output
		.I0(Q_out1426) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1428(
		.O(Q_out1428), // LUT general output
		.I0(Q_out1427) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1429(
		.O(Q_out1429), // LUT general output
		.I0(Q_out1428) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1430(
		.O(Q_out1430), // LUT general output
		.I0(Q_out1429) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1431(
		.O(Q_out1431), // LUT general output
		.I0(Q_out1430) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1432(
		.O(Q_out1432), // LUT general output
		.I0(Q_out1431) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1433(
		.O(Q_out1433), // LUT general output
		.I0(Q_out1432) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1434(
		.O(Q_out1434), // LUT general output
		.I0(Q_out1433) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1435(
		.O(Q_out1435), // LUT general output
		.I0(Q_out1434) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1436(
		.O(Q_out1436), // LUT general output
		.I0(Q_out1435) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1437(
		.O(Q_out1437), // LUT general output
		.I0(Q_out1436) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1438(
		.O(Q_out1438), // LUT general output
		.I0(Q_out1437) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1439(
		.O(Q_out1439), // LUT general output
		.I0(Q_out1438) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1440(
		.O(Q_out1440), // LUT general output
		.I0(Q_out1439) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1441(
		.O(Q_out1441), // LUT general output
		.I0(Q_out1440) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1442(
		.O(Q_out1442), // LUT general output
		.I0(Q_out1441) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1443(
		.O(Q_out1443), // LUT general output
		.I0(Q_out1442) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1444(
		.O(Q_out1444), // LUT general output
		.I0(Q_out1443) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1445(
		.O(Q_out1445), // LUT general output
		.I0(Q_out1444) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1446(
		.O(Q_out1446), // LUT general output
		.I0(Q_out1445) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1447(
		.O(Q_out1447), // LUT general output
		.I0(Q_out1446) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1448(
		.O(Q_out1448), // LUT general output
		.I0(Q_out1447) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1449(
		.O(Q_out1449), // LUT general output
		.I0(Q_out1448) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1450(
		.O(Q_out1450), // LUT general output
		.I0(Q_out1449) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1451(
		.O(Q_out1451), // LUT general output
		.I0(Q_out1450) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1452(
		.O(Q_out1452), // LUT general output
		.I0(Q_out1451) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1453(
		.O(Q_out1453), // LUT general output
		.I0(Q_out1452) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1454(
		.O(Q_out1454), // LUT general output
		.I0(Q_out1453) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1455(
		.O(Q_out1455), // LUT general output
		.I0(Q_out1454) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1456(
		.O(Q_out1456), // LUT general output
		.I0(Q_out1455) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1457(
		.O(Q_out1457), // LUT general output
		.I0(Q_out1456) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1458(
		.O(Q_out1458), // LUT general output
		.I0(Q_out1457) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1459(
		.O(Q_out1459), // LUT general output
		.I0(Q_out1458) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1460(
		.O(Q_out1460), // LUT general output
		.I0(Q_out1459) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1461(
		.O(Q_out1461), // LUT general output
		.I0(Q_out1460) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1462(
		.O(Q_out1462), // LUT general output
		.I0(Q_out1461) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1463(
		.O(Q_out1463), // LUT general output
		.I0(Q_out1462) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1464(
		.O(Q_out1464), // LUT general output
		.I0(Q_out1463) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1465(
		.O(Q_out1465), // LUT general output
		.I0(Q_out1464) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1466(
		.O(Q_out1466), // LUT general output
		.I0(Q_out1465) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1467(
		.O(Q_out1467), // LUT general output
		.I0(Q_out1466) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1468(
		.O(Q_out1468), // LUT general output
		.I0(Q_out1467) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1469(
		.O(Q_out1469), // LUT general output
		.I0(Q_out1468) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1470(
		.O(Q_out1470), // LUT general output
		.I0(Q_out1469) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1471(
		.O(Q_out1471), // LUT general output
		.I0(Q_out1470) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1472(
		.O(Q_out1472), // LUT general output
		.I0(Q_out1471) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1473(
		.O(Q_out1473), // LUT general output
		.I0(Q_out1472) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1474(
		.O(Q_out1474), // LUT general output
		.I0(Q_out1473) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1475(
		.O(Q_out1475), // LUT general output
		.I0(Q_out1474) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1476(
		.O(Q_out1476), // LUT general output
		.I0(Q_out1475) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1477(
		.O(Q_out1477), // LUT general output
		.I0(Q_out1476) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1478(
		.O(Q_out1478), // LUT general output
		.I0(Q_out1477) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1479(
		.O(Q_out1479), // LUT general output
		.I0(Q_out1478) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1480(
		.O(Q_out1480), // LUT general output
		.I0(Q_out1479) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1481(
		.O(Q_out1481), // LUT general output
		.I0(Q_out1480) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1482(
		.O(Q_out1482), // LUT general output
		.I0(Q_out1481) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1483(
		.O(Q_out1483), // LUT general output
		.I0(Q_out1482) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1484(
		.O(Q_out1484), // LUT general output
		.I0(Q_out1483) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1485(
		.O(Q_out1485), // LUT general output
		.I0(Q_out1484) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1486(
		.O(Q_out1486), // LUT general output
		.I0(Q_out1485) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1487(
		.O(Q_out1487), // LUT general output
		.I0(Q_out1486) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1488(
		.O(Q_out1488), // LUT general output
		.I0(Q_out1487) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1489(
		.O(Q_out1489), // LUT general output
		.I0(Q_out1488) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1490(
		.O(Q_out1490), // LUT general output
		.I0(Q_out1489) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1491(
		.O(Q_out1491), // LUT general output
		.I0(Q_out1490) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1492(
		.O(Q_out1492), // LUT general output
		.I0(Q_out1491) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1493(
		.O(Q_out1493), // LUT general output
		.I0(Q_out1492) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1494(
		.O(Q_out1494), // LUT general output
		.I0(Q_out1493) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1495(
		.O(Q_out1495), // LUT general output
		.I0(Q_out1494) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1496(
		.O(Q_out1496), // LUT general output
		.I0(Q_out1495) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1497(
		.O(Q_out1497), // LUT general output
		.I0(Q_out1496) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1498(
		.O(Q_out1498), // LUT general output
		.I0(Q_out1497) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1499(
		.O(Q_out1499), // LUT general output
		.I0(Q_out1498) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1500(
		.O(Q_out1500), // LUT general output
		.I0(Q_out1499) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1501(
		.O(Q_out1501), // LUT general output
		.I0(Q_out1500) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1502(
		.O(Q_out1502), // LUT general output
		.I0(Q_out1501) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1503(
		.O(Q_out1503), // LUT general output
		.I0(Q_out1502) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1504(
		.O(Q_out1504), // LUT general output
		.I0(Q_out1503) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1505(
		.O(Q_out1505), // LUT general output
		.I0(Q_out1504) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1506(
		.O(Q_out1506), // LUT general output
		.I0(Q_out1505) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1507(
		.O(Q_out1507), // LUT general output
		.I0(Q_out1506) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1508(
		.O(Q_out1508), // LUT general output
		.I0(Q_out1507) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1509(
		.O(Q_out1509), // LUT general output
		.I0(Q_out1508) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1510(
		.O(Q_out1510), // LUT general output
		.I0(Q_out1509) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1511(
		.O(Q_out1511), // LUT general output
		.I0(Q_out1510) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1512(
		.O(Q_out1512), // LUT general output
		.I0(Q_out1511) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1513(
		.O(Q_out1513), // LUT general output
		.I0(Q_out1512) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1514(
		.O(Q_out1514), // LUT general output
		.I0(Q_out1513) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1515(
		.O(Q_out1515), // LUT general output
		.I0(Q_out1514) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1516(
		.O(Q_out1516), // LUT general output
		.I0(Q_out1515) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1517(
		.O(Q_out1517), // LUT general output
		.I0(Q_out1516) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1518(
		.O(Q_out1518), // LUT general output
		.I0(Q_out1517) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1519(
		.O(Q_out1519), // LUT general output
		.I0(Q_out1518) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1520(
		.O(Q_out1520), // LUT general output
		.I0(Q_out1519) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1521(
		.O(Q_out1521), // LUT general output
		.I0(Q_out1520) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1522(
		.O(Q_out1522), // LUT general output
		.I0(Q_out1521) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1523(
		.O(Q_out1523), // LUT general output
		.I0(Q_out1522) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1524(
		.O(Q_out1524), // LUT general output
		.I0(Q_out1523) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1525(
		.O(Q_out1525), // LUT general output
		.I0(Q_out1524) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1526(
		.O(Q_out1526), // LUT general output
		.I0(Q_out1525) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1527(
		.O(Q_out1527), // LUT general output
		.I0(Q_out1526) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1528(
		.O(Q_out1528), // LUT general output
		.I0(Q_out1527) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1529(
		.O(Q_out1529), // LUT general output
		.I0(Q_out1528) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1530(
		.O(Q_out1530), // LUT general output
		.I0(Q_out1529) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1531(
		.O(Q_out1531), // LUT general output
		.I0(Q_out1530) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1532(
		.O(Q_out1532), // LUT general output
		.I0(Q_out1531) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1533(
		.O(Q_out1533), // LUT general output
		.I0(Q_out1532) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1534(
		.O(Q_out1534), // LUT general output
		.I0(Q_out1533) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1535(
		.O(Q_out1535), // LUT general output
		.I0(Q_out1534) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1536(
		.O(Q_out1536), // LUT general output
		.I0(Q_out1535) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1537(
		.O(Q_out1537), // LUT general output
		.I0(Q_out1536) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1538(
		.O(Q_out1538), // LUT general output
		.I0(Q_out1537) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1539(
		.O(Q_out1539), // LUT general output
		.I0(Q_out1538) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1540(
		.O(Q_out1540), // LUT general output
		.I0(Q_out1539) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1541(
		.O(Q_out1541), // LUT general output
		.I0(Q_out1540) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1542(
		.O(Q_out1542), // LUT general output
		.I0(Q_out1541) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1543(
		.O(Q_out1543), // LUT general output
		.I0(Q_out1542) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1544(
		.O(Q_out1544), // LUT general output
		.I0(Q_out1543) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1545(
		.O(Q_out1545), // LUT general output
		.I0(Q_out1544) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1546(
		.O(Q_out1546), // LUT general output
		.I0(Q_out1545) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1547(
		.O(Q_out1547), // LUT general output
		.I0(Q_out1546) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1548(
		.O(Q_out1548), // LUT general output
		.I0(Q_out1547) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1549(
		.O(Q_out1549), // LUT general output
		.I0(Q_out1548) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1550(
		.O(Q_out1550), // LUT general output
		.I0(Q_out1549) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1551(
		.O(Q_out1551), // LUT general output
		.I0(Q_out1550) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1552(
		.O(Q_out1552), // LUT general output
		.I0(Q_out1551) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1553(
		.O(Q_out1553), // LUT general output
		.I0(Q_out1552) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1554(
		.O(Q_out1554), // LUT general output
		.I0(Q_out1553) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1555(
		.O(Q_out1555), // LUT general output
		.I0(Q_out1554) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1556(
		.O(Q_out1556), // LUT general output
		.I0(Q_out1555) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1557(
		.O(Q_out1557), // LUT general output
		.I0(Q_out1556) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1558(
		.O(Q_out1558), // LUT general output
		.I0(Q_out1557) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1559(
		.O(Q_out1559), // LUT general output
		.I0(Q_out1558) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1560(
		.O(Q_out1560), // LUT general output
		.I0(Q_out1559) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1561(
		.O(Q_out1561), // LUT general output
		.I0(Q_out1560) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1562(
		.O(Q_out1562), // LUT general output
		.I0(Q_out1561) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1563(
		.O(Q_out1563), // LUT general output
		.I0(Q_out1562) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1564(
		.O(Q_out1564), // LUT general output
		.I0(Q_out1563) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1565(
		.O(Q_out1565), // LUT general output
		.I0(Q_out1564) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1566(
		.O(Q_out1566), // LUT general output
		.I0(Q_out1565) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1567(
		.O(Q_out1567), // LUT general output
		.I0(Q_out1566) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1568(
		.O(Q_out1568), // LUT general output
		.I0(Q_out1567) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1569(
		.O(Q_out1569), // LUT general output
		.I0(Q_out1568) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1570(
		.O(Q_out1570), // LUT general output
		.I0(Q_out1569) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1571(
		.O(Q_out1571), // LUT general output
		.I0(Q_out1570) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1572(
		.O(Q_out1572), // LUT general output
		.I0(Q_out1571) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1573(
		.O(Q_out1573), // LUT general output
		.I0(Q_out1572) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1574(
		.O(Q_out1574), // LUT general output
		.I0(Q_out1573) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1575(
		.O(Q_out1575), // LUT general output
		.I0(Q_out1574) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1576(
		.O(Q_out1576), // LUT general output
		.I0(Q_out1575) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1577(
		.O(Q_out1577), // LUT general output
		.I0(Q_out1576) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1578(
		.O(Q_out1578), // LUT general output
		.I0(Q_out1577) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1579(
		.O(Q_out1579), // LUT general output
		.I0(Q_out1578) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1580(
		.O(Q_out1580), // LUT general output
		.I0(Q_out1579) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1581(
		.O(Q_out1581), // LUT general output
		.I0(Q_out1580) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1582(
		.O(Q_out1582), // LUT general output
		.I0(Q_out1581) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1583(
		.O(Q_out1583), // LUT general output
		.I0(Q_out1582) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1584(
		.O(Q_out1584), // LUT general output
		.I0(Q_out1583) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1585(
		.O(Q_out1585), // LUT general output
		.I0(Q_out1584) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1586(
		.O(Q_out1586), // LUT general output
		.I0(Q_out1585) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1587(
		.O(Q_out1587), // LUT general output
		.I0(Q_out1586) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1588(
		.O(Q_out1588), // LUT general output
		.I0(Q_out1587) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1589(
		.O(Q_out1589), // LUT general output
		.I0(Q_out1588) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1590(
		.O(Q_out1590), // LUT general output
		.I0(Q_out1589) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1591(
		.O(Q_out1591), // LUT general output
		.I0(Q_out1590) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1592(
		.O(Q_out1592), // LUT general output
		.I0(Q_out1591) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1593(
		.O(Q_out1593), // LUT general output
		.I0(Q_out1592) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1594(
		.O(Q_out1594), // LUT general output
		.I0(Q_out1593) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1595(
		.O(Q_out1595), // LUT general output
		.I0(Q_out1594) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1596(
		.O(Q_out1596), // LUT general output
		.I0(Q_out1595) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1597(
		.O(Q_out1597), // LUT general output
		.I0(Q_out1596) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1598(
		.O(Q_out1598), // LUT general output
		.I0(Q_out1597) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1599(
		.O(Q_out1599), // LUT general output
		.I0(Q_out1598) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1600(
		.O(Q_out1600), // LUT general output
		.I0(Q_out1599) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1601(
		.O(Q_out1601), // LUT general output
		.I0(Q_out1600) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1602(
		.O(Q_out1602), // LUT general output
		.I0(Q_out1601) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1603(
		.O(Q_out1603), // LUT general output
		.I0(Q_out1602) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1604(
		.O(Q_out1604), // LUT general output
		.I0(Q_out1603) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1605(
		.O(Q_out1605), // LUT general output
		.I0(Q_out1604) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1606(
		.O(Q_out1606), // LUT general output
		.I0(Q_out1605) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1607(
		.O(Q_out1607), // LUT general output
		.I0(Q_out1606) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1608(
		.O(Q_out1608), // LUT general output
		.I0(Q_out1607) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1609(
		.O(Q_out1609), // LUT general output
		.I0(Q_out1608) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1610(
		.O(Q_out1610), // LUT general output
		.I0(Q_out1609) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1611(
		.O(Q_out1611), // LUT general output
		.I0(Q_out1610) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1612(
		.O(Q_out1612), // LUT general output
		.I0(Q_out1611) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1613(
		.O(Q_out1613), // LUT general output
		.I0(Q_out1612) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1614(
		.O(Q_out1614), // LUT general output
		.I0(Q_out1613) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1615(
		.O(Q_out1615), // LUT general output
		.I0(Q_out1614) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1616(
		.O(Q_out1616), // LUT general output
		.I0(Q_out1615) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1617(
		.O(Q_out1617), // LUT general output
		.I0(Q_out1616) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1618(
		.O(Q_out1618), // LUT general output
		.I0(Q_out1617) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1619(
		.O(Q_out1619), // LUT general output
		.I0(Q_out1618) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1620(
		.O(Q_out1620), // LUT general output
		.I0(Q_out1619) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1621(
		.O(Q_out1621), // LUT general output
		.I0(Q_out1620) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1622(
		.O(Q_out1622), // LUT general output
		.I0(Q_out1621) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1623(
		.O(Q_out1623), // LUT general output
		.I0(Q_out1622) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1624(
		.O(Q_out1624), // LUT general output
		.I0(Q_out1623) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1625(
		.O(Q_out1625), // LUT general output
		.I0(Q_out1624) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1626(
		.O(Q_out1626), // LUT general output
		.I0(Q_out1625) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1627(
		.O(Q_out1627), // LUT general output
		.I0(Q_out1626) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1628(
		.O(Q_out1628), // LUT general output
		.I0(Q_out1627) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1629(
		.O(Q_out1629), // LUT general output
		.I0(Q_out1628) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1630(
		.O(Q_out1630), // LUT general output
		.I0(Q_out1629) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1631(
		.O(Q_out1631), // LUT general output
		.I0(Q_out1630) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1632(
		.O(Q_out1632), // LUT general output
		.I0(Q_out1631) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1633(
		.O(Q_out1633), // LUT general output
		.I0(Q_out1632) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1634(
		.O(Q_out1634), // LUT general output
		.I0(Q_out1633) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1635(
		.O(Q_out1635), // LUT general output
		.I0(Q_out1634) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1636(
		.O(Q_out1636), // LUT general output
		.I0(Q_out1635) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1637(
		.O(Q_out1637), // LUT general output
		.I0(Q_out1636) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1638(
		.O(Q_out1638), // LUT general output
		.I0(Q_out1637) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1639(
		.O(Q_out1639), // LUT general output
		.I0(Q_out1638) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1640(
		.O(Q_out1640), // LUT general output
		.I0(Q_out1639) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1641(
		.O(Q_out1641), // LUT general output
		.I0(Q_out1640) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1642(
		.O(Q_out1642), // LUT general output
		.I0(Q_out1641) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1643(
		.O(Q_out1643), // LUT general output
		.I0(Q_out1642) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1644(
		.O(Q_out1644), // LUT general output
		.I0(Q_out1643) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1645(
		.O(Q_out1645), // LUT general output
		.I0(Q_out1644) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1646(
		.O(Q_out1646), // LUT general output
		.I0(Q_out1645) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1647(
		.O(Q_out1647), // LUT general output
		.I0(Q_out1646) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1648(
		.O(Q_out1648), // LUT general output
		.I0(Q_out1647) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1649(
		.O(Q_out1649), // LUT general output
		.I0(Q_out1648) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1650(
		.O(Q_out1650), // LUT general output
		.I0(Q_out1649) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1651(
		.O(Q_out1651), // LUT general output
		.I0(Q_out1650) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1652(
		.O(Q_out1652), // LUT general output
		.I0(Q_out1651) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1653(
		.O(Q_out1653), // LUT general output
		.I0(Q_out1652) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1654(
		.O(Q_out1654), // LUT general output
		.I0(Q_out1653) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1655(
		.O(Q_out1655), // LUT general output
		.I0(Q_out1654) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1656(
		.O(Q_out1656), // LUT general output
		.I0(Q_out1655) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1657(
		.O(Q_out1657), // LUT general output
		.I0(Q_out1656) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1658(
		.O(Q_out1658), // LUT general output
		.I0(Q_out1657) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1659(
		.O(Q_out1659), // LUT general output
		.I0(Q_out1658) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1660(
		.O(Q_out1660), // LUT general output
		.I0(Q_out1659) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1661(
		.O(Q_out1661), // LUT general output
		.I0(Q_out1660) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1662(
		.O(Q_out1662), // LUT general output
		.I0(Q_out1661) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1663(
		.O(Q_out1663), // LUT general output
		.I0(Q_out1662) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1664(
		.O(Q_out1664), // LUT general output
		.I0(Q_out1663) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1665(
		.O(Q_out1665), // LUT general output
		.I0(Q_out1664) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1666(
		.O(Q_out1666), // LUT general output
		.I0(Q_out1665) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1667(
		.O(Q_out1667), // LUT general output
		.I0(Q_out1666) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1668(
		.O(Q_out1668), // LUT general output
		.I0(Q_out1667) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1669(
		.O(Q_out1669), // LUT general output
		.I0(Q_out1668) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1670(
		.O(Q_out1670), // LUT general output
		.I0(Q_out1669) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1671(
		.O(Q_out1671), // LUT general output
		.I0(Q_out1670) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1672(
		.O(Q_out1672), // LUT general output
		.I0(Q_out1671) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1673(
		.O(Q_out1673), // LUT general output
		.I0(Q_out1672) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1674(
		.O(Q_out1674), // LUT general output
		.I0(Q_out1673) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1675(
		.O(Q_out1675), // LUT general output
		.I0(Q_out1674) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1676(
		.O(Q_out1676), // LUT general output
		.I0(Q_out1675) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1677(
		.O(Q_out1677), // LUT general output
		.I0(Q_out1676) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1678(
		.O(Q_out1678), // LUT general output
		.I0(Q_out1677) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1679(
		.O(Q_out1679), // LUT general output
		.I0(Q_out1678) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1680(
		.O(Q_out1680), // LUT general output
		.I0(Q_out1679) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1681(
		.O(Q_out1681), // LUT general output
		.I0(Q_out1680) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1682(
		.O(Q_out1682), // LUT general output
		.I0(Q_out1681) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1683(
		.O(Q_out1683), // LUT general output
		.I0(Q_out1682) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1684(
		.O(Q_out1684), // LUT general output
		.I0(Q_out1683) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1685(
		.O(Q_out1685), // LUT general output
		.I0(Q_out1684) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1686(
		.O(Q_out1686), // LUT general output
		.I0(Q_out1685) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1687(
		.O(Q_out1687), // LUT general output
		.I0(Q_out1686) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1688(
		.O(Q_out1688), // LUT general output
		.I0(Q_out1687) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1689(
		.O(Q_out1689), // LUT general output
		.I0(Q_out1688) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1690(
		.O(Q_out1690), // LUT general output
		.I0(Q_out1689) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1691(
		.O(Q_out1691), // LUT general output
		.I0(Q_out1690) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1692(
		.O(Q_out1692), // LUT general output
		.I0(Q_out1691) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1693(
		.O(Q_out1693), // LUT general output
		.I0(Q_out1692) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1694(
		.O(Q_out1694), // LUT general output
		.I0(Q_out1693) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1695(
		.O(Q_out1695), // LUT general output
		.I0(Q_out1694) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1696(
		.O(Q_out1696), // LUT general output
		.I0(Q_out1695) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1697(
		.O(Q_out1697), // LUT general output
		.I0(Q_out1696) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1698(
		.O(Q_out1698), // LUT general output
		.I0(Q_out1697) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1699(
		.O(Q_out1699), // LUT general output
		.I0(Q_out1698) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1700(
		.O(Q_out1700), // LUT general output
		.I0(Q_out1699) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1701(
		.O(Q_out1701), // LUT general output
		.I0(Q_out1700) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1702(
		.O(Q_out1702), // LUT general output
		.I0(Q_out1701) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1703(
		.O(Q_out1703), // LUT general output
		.I0(Q_out1702) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1704(
		.O(Q_out1704), // LUT general output
		.I0(Q_out1703) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1705(
		.O(Q_out1705), // LUT general output
		.I0(Q_out1704) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1706(
		.O(Q_out1706), // LUT general output
		.I0(Q_out1705) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1707(
		.O(Q_out1707), // LUT general output
		.I0(Q_out1706) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1708(
		.O(Q_out1708), // LUT general output
		.I0(Q_out1707) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1709(
		.O(Q_out1709), // LUT general output
		.I0(Q_out1708) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1710(
		.O(Q_out1710), // LUT general output
		.I0(Q_out1709) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1711(
		.O(Q_out1711), // LUT general output
		.I0(Q_out1710) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1712(
		.O(Q_out1712), // LUT general output
		.I0(Q_out1711) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1713(
		.O(Q_out1713), // LUT general output
		.I0(Q_out1712) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1714(
		.O(Q_out1714), // LUT general output
		.I0(Q_out1713) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1715(
		.O(Q_out1715), // LUT general output
		.I0(Q_out1714) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1716(
		.O(Q_out1716), // LUT general output
		.I0(Q_out1715) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1717(
		.O(Q_out1717), // LUT general output
		.I0(Q_out1716) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1718(
		.O(Q_out1718), // LUT general output
		.I0(Q_out1717) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1719(
		.O(Q_out1719), // LUT general output
		.I0(Q_out1718) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1720(
		.O(Q_out1720), // LUT general output
		.I0(Q_out1719) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1721(
		.O(Q_out1721), // LUT general output
		.I0(Q_out1720) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1722(
		.O(Q_out1722), // LUT general output
		.I0(Q_out1721) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1723(
		.O(Q_out1723), // LUT general output
		.I0(Q_out1722) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1724(
		.O(Q_out1724), // LUT general output
		.I0(Q_out1723) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1725(
		.O(Q_out1725), // LUT general output
		.I0(Q_out1724) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1726(
		.O(Q_out1726), // LUT general output
		.I0(Q_out1725) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1727(
		.O(Q_out1727), // LUT general output
		.I0(Q_out1726) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1728(
		.O(Q_out1728), // LUT general output
		.I0(Q_out1727) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1729(
		.O(Q_out1729), // LUT general output
		.I0(Q_out1728) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1730(
		.O(Q_out1730), // LUT general output
		.I0(Q_out1729) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1731(
		.O(Q_out1731), // LUT general output
		.I0(Q_out1730) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1732(
		.O(Q_out1732), // LUT general output
		.I0(Q_out1731) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1733(
		.O(Q_out1733), // LUT general output
		.I0(Q_out1732) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1734(
		.O(Q_out1734), // LUT general output
		.I0(Q_out1733) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1735(
		.O(Q_out1735), // LUT general output
		.I0(Q_out1734) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1736(
		.O(Q_out1736), // LUT general output
		.I0(Q_out1735) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1737(
		.O(Q_out1737), // LUT general output
		.I0(Q_out1736) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1738(
		.O(Q_out1738), // LUT general output
		.I0(Q_out1737) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1739(
		.O(Q_out1739), // LUT general output
		.I0(Q_out1738) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1740(
		.O(Q_out1740), // LUT general output
		.I0(Q_out1739) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1741(
		.O(Q_out1741), // LUT general output
		.I0(Q_out1740) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1742(
		.O(Q_out1742), // LUT general output
		.I0(Q_out1741) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1743(
		.O(Q_out1743), // LUT general output
		.I0(Q_out1742) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1744(
		.O(Q_out1744), // LUT general output
		.I0(Q_out1743) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1745(
		.O(Q_out1745), // LUT general output
		.I0(Q_out1744) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1746(
		.O(Q_out1746), // LUT general output
		.I0(Q_out1745) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1747(
		.O(Q_out1747), // LUT general output
		.I0(Q_out1746) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1748(
		.O(Q_out1748), // LUT general output
		.I0(Q_out1747) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1749(
		.O(Q_out1749), // LUT general output
		.I0(Q_out1748) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1750(
		.O(Q_out1750), // LUT general output
		.I0(Q_out1749) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1751(
		.O(Q_out1751), // LUT general output
		.I0(Q_out1750) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1752(
		.O(Q_out1752), // LUT general output
		.I0(Q_out1751) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1753(
		.O(Q_out1753), // LUT general output
		.I0(Q_out1752) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1754(
		.O(Q_out1754), // LUT general output
		.I0(Q_out1753) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1755(
		.O(Q_out1755), // LUT general output
		.I0(Q_out1754) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1756(
		.O(Q_out1756), // LUT general output
		.I0(Q_out1755) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1757(
		.O(Q_out1757), // LUT general output
		.I0(Q_out1756) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1758(
		.O(Q_out1758), // LUT general output
		.I0(Q_out1757) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1759(
		.O(Q_out1759), // LUT general output
		.I0(Q_out1758) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1760(
		.O(Q_out1760), // LUT general output
		.I0(Q_out1759) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1761(
		.O(Q_out1761), // LUT general output
		.I0(Q_out1760) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1762(
		.O(Q_out1762), // LUT general output
		.I0(Q_out1761) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1763(
		.O(Q_out1763), // LUT general output
		.I0(Q_out1762) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1764(
		.O(Q_out1764), // LUT general output
		.I0(Q_out1763) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1765(
		.O(Q_out1765), // LUT general output
		.I0(Q_out1764) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1766(
		.O(Q_out1766), // LUT general output
		.I0(Q_out1765) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1767(
		.O(Q_out1767), // LUT general output
		.I0(Q_out1766) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1768(
		.O(Q_out1768), // LUT general output
		.I0(Q_out1767) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1769(
		.O(Q_out1769), // LUT general output
		.I0(Q_out1768) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1770(
		.O(Q_out1770), // LUT general output
		.I0(Q_out1769) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1771(
		.O(Q_out1771), // LUT general output
		.I0(Q_out1770) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1772(
		.O(Q_out1772), // LUT general output
		.I0(Q_out1771) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1773(
		.O(Q_out1773), // LUT general output
		.I0(Q_out1772) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1774(
		.O(Q_out1774), // LUT general output
		.I0(Q_out1773) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1775(
		.O(Q_out1775), // LUT general output
		.I0(Q_out1774) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1776(
		.O(Q_out1776), // LUT general output
		.I0(Q_out1775) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1777(
		.O(Q_out1777), // LUT general output
		.I0(Q_out1776) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1778(
		.O(Q_out1778), // LUT general output
		.I0(Q_out1777) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1779(
		.O(Q_out1779), // LUT general output
		.I0(Q_out1778) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1780(
		.O(Q_out1780), // LUT general output
		.I0(Q_out1779) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1781(
		.O(Q_out1781), // LUT general output
		.I0(Q_out1780) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1782(
		.O(Q_out1782), // LUT general output
		.I0(Q_out1781) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1783(
		.O(Q_out1783), // LUT general output
		.I0(Q_out1782) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1784(
		.O(Q_out1784), // LUT general output
		.I0(Q_out1783) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1785(
		.O(Q_out1785), // LUT general output
		.I0(Q_out1784) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1786(
		.O(Q_out1786), // LUT general output
		.I0(Q_out1785) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1787(
		.O(Q_out1787), // LUT general output
		.I0(Q_out1786) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1788(
		.O(Q_out1788), // LUT general output
		.I0(Q_out1787) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1789(
		.O(Q_out1789), // LUT general output
		.I0(Q_out1788) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1790(
		.O(Q_out1790), // LUT general output
		.I0(Q_out1789) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1791(
		.O(Q_out1791), // LUT general output
		.I0(Q_out1790) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1792(
		.O(Q_out1792), // LUT general output
		.I0(Q_out1791) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1793(
		.O(Q_out1793), // LUT general output
		.I0(Q_out1792) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1794(
		.O(Q_out1794), // LUT general output
		.I0(Q_out1793) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1795(
		.O(Q_out1795), // LUT general output
		.I0(Q_out1794) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1796(
		.O(Q_out1796), // LUT general output
		.I0(Q_out1795) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1797(
		.O(Q_out1797), // LUT general output
		.I0(Q_out1796) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1798(
		.O(Q_out1798), // LUT general output
		.I0(Q_out1797) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1799(
		.O(Q_out1799), // LUT general output
		.I0(Q_out1798) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1800(
		.O(Q_out1800), // LUT general output
		.I0(Q_out1799) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1801(
		.O(Q_out1801), // LUT general output
		.I0(Q_out1800) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1802(
		.O(Q_out1802), // LUT general output
		.I0(Q_out1801) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1803(
		.O(Q_out1803), // LUT general output
		.I0(Q_out1802) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1804(
		.O(Q_out1804), // LUT general output
		.I0(Q_out1803) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1805(
		.O(Q_out1805), // LUT general output
		.I0(Q_out1804) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1806(
		.O(Q_out1806), // LUT general output
		.I0(Q_out1805) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1807(
		.O(Q_out1807), // LUT general output
		.I0(Q_out1806) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1808(
		.O(Q_out1808), // LUT general output
		.I0(Q_out1807) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1809(
		.O(Q_out1809), // LUT general output
		.I0(Q_out1808) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1810(
		.O(Q_out1810), // LUT general output
		.I0(Q_out1809) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1811(
		.O(Q_out1811), // LUT general output
		.I0(Q_out1810) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1812(
		.O(Q_out1812), // LUT general output
		.I0(Q_out1811) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1813(
		.O(Q_out1813), // LUT general output
		.I0(Q_out1812) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1814(
		.O(Q_out1814), // LUT general output
		.I0(Q_out1813) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1815(
		.O(Q_out1815), // LUT general output
		.I0(Q_out1814) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1816(
		.O(Q_out1816), // LUT general output
		.I0(Q_out1815) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1817(
		.O(Q_out1817), // LUT general output
		.I0(Q_out1816) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1818(
		.O(Q_out1818), // LUT general output
		.I0(Q_out1817) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1819(
		.O(Q_out1819), // LUT general output
		.I0(Q_out1818) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1820(
		.O(Q_out1820), // LUT general output
		.I0(Q_out1819) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1821(
		.O(Q_out1821), // LUT general output
		.I0(Q_out1820) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1822(
		.O(Q_out1822), // LUT general output
		.I0(Q_out1821) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1823(
		.O(Q_out1823), // LUT general output
		.I0(Q_out1822) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1824(
		.O(Q_out1824), // LUT general output
		.I0(Q_out1823) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1825(
		.O(Q_out1825), // LUT general output
		.I0(Q_out1824) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1826(
		.O(Q_out1826), // LUT general output
		.I0(Q_out1825) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1827(
		.O(Q_out1827), // LUT general output
		.I0(Q_out1826) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1828(
		.O(Q_out1828), // LUT general output
		.I0(Q_out1827) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1829(
		.O(Q_out1829), // LUT general output
		.I0(Q_out1828) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1830(
		.O(Q_out1830), // LUT general output
		.I0(Q_out1829) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1831(
		.O(Q_out1831), // LUT general output
		.I0(Q_out1830) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1832(
		.O(Q_out1832), // LUT general output
		.I0(Q_out1831) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1833(
		.O(Q_out1833), // LUT general output
		.I0(Q_out1832) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1834(
		.O(Q_out1834), // LUT general output
		.I0(Q_out1833) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1835(
		.O(Q_out1835), // LUT general output
		.I0(Q_out1834) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1836(
		.O(Q_out1836), // LUT general output
		.I0(Q_out1835) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1837(
		.O(Q_out1837), // LUT general output
		.I0(Q_out1836) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1838(
		.O(Q_out1838), // LUT general output
		.I0(Q_out1837) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1839(
		.O(Q_out1839), // LUT general output
		.I0(Q_out1838) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1840(
		.O(Q_out1840), // LUT general output
		.I0(Q_out1839) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1841(
		.O(Q_out1841), // LUT general output
		.I0(Q_out1840) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1842(
		.O(Q_out1842), // LUT general output
		.I0(Q_out1841) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1843(
		.O(Q_out1843), // LUT general output
		.I0(Q_out1842) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1844(
		.O(Q_out1844), // LUT general output
		.I0(Q_out1843) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1845(
		.O(Q_out1845), // LUT general output
		.I0(Q_out1844) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1846(
		.O(Q_out1846), // LUT general output
		.I0(Q_out1845) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1847(
		.O(Q_out1847), // LUT general output
		.I0(Q_out1846) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1848(
		.O(Q_out1848), // LUT general output
		.I0(Q_out1847) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1849(
		.O(Q_out1849), // LUT general output
		.I0(Q_out1848) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1850(
		.O(Q_out1850), // LUT general output
		.I0(Q_out1849) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1851(
		.O(Q_out1851), // LUT general output
		.I0(Q_out1850) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1852(
		.O(Q_out1852), // LUT general output
		.I0(Q_out1851) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1853(
		.O(Q_out1853), // LUT general output
		.I0(Q_out1852) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1854(
		.O(Q_out1854), // LUT general output
		.I0(Q_out1853) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1855(
		.O(Q_out1855), // LUT general output
		.I0(Q_out1854) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1856(
		.O(Q_out1856), // LUT general output
		.I0(Q_out1855) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1857(
		.O(Q_out1857), // LUT general output
		.I0(Q_out1856) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1858(
		.O(Q_out1858), // LUT general output
		.I0(Q_out1857) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1859(
		.O(Q_out1859), // LUT general output
		.I0(Q_out1858) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1860(
		.O(Q_out1860), // LUT general output
		.I0(Q_out1859) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1861(
		.O(Q_out1861), // LUT general output
		.I0(Q_out1860) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1862(
		.O(Q_out1862), // LUT general output
		.I0(Q_out1861) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1863(
		.O(Q_out1863), // LUT general output
		.I0(Q_out1862) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1864(
		.O(Q_out1864), // LUT general output
		.I0(Q_out1863) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1865(
		.O(Q_out1865), // LUT general output
		.I0(Q_out1864) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1866(
		.O(Q_out1866), // LUT general output
		.I0(Q_out1865) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1867(
		.O(Q_out1867), // LUT general output
		.I0(Q_out1866) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1868(
		.O(Q_out1868), // LUT general output
		.I0(Q_out1867) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1869(
		.O(Q_out1869), // LUT general output
		.I0(Q_out1868) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1870(
		.O(Q_out1870), // LUT general output
		.I0(Q_out1869) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1871(
		.O(Q_out1871), // LUT general output
		.I0(Q_out1870) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1872(
		.O(Q_out1872), // LUT general output
		.I0(Q_out1871) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1873(
		.O(Q_out1873), // LUT general output
		.I0(Q_out1872) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1874(
		.O(Q_out1874), // LUT general output
		.I0(Q_out1873) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1875(
		.O(Q_out1875), // LUT general output
		.I0(Q_out1874) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1876(
		.O(Q_out1876), // LUT general output
		.I0(Q_out1875) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1877(
		.O(Q_out1877), // LUT general output
		.I0(Q_out1876) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1878(
		.O(Q_out1878), // LUT general output
		.I0(Q_out1877) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1879(
		.O(Q_out1879), // LUT general output
		.I0(Q_out1878) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1880(
		.O(Q_out1880), // LUT general output
		.I0(Q_out1879) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1881(
		.O(Q_out1881), // LUT general output
		.I0(Q_out1880) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1882(
		.O(Q_out1882), // LUT general output
		.I0(Q_out1881) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1883(
		.O(Q_out1883), // LUT general output
		.I0(Q_out1882) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1884(
		.O(Q_out1884), // LUT general output
		.I0(Q_out1883) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1885(
		.O(Q_out1885), // LUT general output
		.I0(Q_out1884) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1886(
		.O(Q_out1886), // LUT general output
		.I0(Q_out1885) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1887(
		.O(Q_out1887), // LUT general output
		.I0(Q_out1886) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1888(
		.O(Q_out1888), // LUT general output
		.I0(Q_out1887) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1889(
		.O(Q_out1889), // LUT general output
		.I0(Q_out1888) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1890(
		.O(Q_out1890), // LUT general output
		.I0(Q_out1889) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1891(
		.O(Q_out1891), // LUT general output
		.I0(Q_out1890) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1892(
		.O(Q_out1892), // LUT general output
		.I0(Q_out1891) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1893(
		.O(Q_out1893), // LUT general output
		.I0(Q_out1892) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1894(
		.O(Q_out1894), // LUT general output
		.I0(Q_out1893) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1895(
		.O(Q_out1895), // LUT general output
		.I0(Q_out1894) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1896(
		.O(Q_out1896), // LUT general output
		.I0(Q_out1895) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1897(
		.O(Q_out1897), // LUT general output
		.I0(Q_out1896) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1898(
		.O(Q_out1898), // LUT general output
		.I0(Q_out1897) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1899(
		.O(Q_out1899), // LUT general output
		.I0(Q_out1898) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_inst1900(
		.O(Q_out1900), // LUT general output
		.I0(Q_out1899) // LUT input
	);


	LUT6 #(
		.INIT(64'h8000000000000001) // BT: this configuration sets O high if all inputs equal
	) LUT6_1 (
		.O(EQUAL), // 1-bit LUT6 output
		.I0(Q_out1), // LUT input
		.I1(Q_out66),  // LUT input
		.I2(Q_out133), // LUT input
		.I3(Q_out200), // LUT input
		.I4(Q_out266), // LUT input
		.I5(Q_out333)  // 1-bit LUT input (fast MUX select only available to O6 output)
	);
		
	LUT6 #(
		.INIT(64'h8000000000000001) 
	) LUT6_2 (
		.O(EQUAL1), // 1-bit LUT6 output
		.I0(Q_out400), // LUT input
		.I1(Q_out466), // LUT input
		.I2(Q_out533), // LUT input
		.I3(Q_out599), // LUT input
		.I4(Q_out666), // LUT input
		.I5(Q_out733)  // 1-bit LUT input (fast MUX select only available to O6 output)
	);
		
	LUT6 #(
		.INIT(64'h8000000000000001) 
	) LUT6_3 (
		.O(EQUAL2), // 1-bit LUT6 output
		.I0(Q_out799),  // LUT input
		.I1(Q_out866),  // LUT input
		.I2(Q_out932),  // LUT input
		.I3(Q_out999),  // LUT input
		.I4(Q_out1066), // LUT input
		.I5(Q_out1132)  // 1-bit LUT input (fast MUX select only available to O6 output)
	);

	
	LUT6 #(
		.INIT(64'h8000000000000001) 
	) LUT6_4 (
		.O(EQUAL3), // 1-bit LUT6 output
		.I0(Q_out1198), // LUT input
		.I1(Q_out1265), // LUT input
		.I2(Q_out1332), // LUT input
		.I3(Q_out1399), // LUT input
		.I4(Q_out1465), // LUT input
		.I5(Q_out1531)  // 1-bit LUT input (fast MUX select only available to O6 output)
	);
		
	LUT6 #(
		.INIT(64'h8000000000000001) 
	) LUT6_5 (
		.O(EQUAL4), // 1-bit LUT6 output
		.I0(Q_out1598), // LUT input
		.I1(Q_out1665), // LUT input
		.I2(Q_out1732), // LUT input
		.I3(Q_out1798), // LUT input
		.I4(Q_out1864), // LUT input
		.I5(Q_out1900)  // 1-bit LUT input (fast MUX select only available to O6 output)
	);
	
	LUT6 #(
		.INIT(64'h8000000000000001) 
	) LUT6_6 (
		.O(CLK_IND), // 1-bit LUT6 output
		.I0(Q_out333),  // LUT input
		.I1(Q_out666),  // LUT input
		.I2(Q_out999),  // LUT input
		.I3(Q_out1333), // LUT input
		.I4(Q_out1666), // LUT input
		.I5(Q_out1900)  // 1-bit LUT input (fast MUX select only available to O6 output)
	);
	
	
	LUT6 #(
		.INIT(64'h8000000000000000) // BT: this configuration sets O high if all inputs high
	) LUT6_7 (
		.O(stop_detect), // 1-bit LUT6 output
		.I0(EQUAL), // LUT input
		.I1(EQUAL1), // LUT input
		.I2(EQUAL2), // LUT input
		.I3(EQUAL3), // LUT input
		.I4(EQUAL4), // LUT input
		.I5(CLK_IND)  // 1-bit LUT input (fast MUX select only available to O6 output)
	);
	

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_dpinst0(
		.O(Q_out_dp0), // LUT general output
		.I0(stop_detect) // LUT input
	);
	
LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_dpinst1(
		.O(Q_out_dp1), // LUT general output
		.I0(Q_out_dp0) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_dpinst2(
		.O(Q_out_dp2), // LUT general output
		.I0(Q_out_dp1) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_dpinst3(
		.O(Q_out_dp3), // LUT general output
		.I0(Q_out_dp2) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_dpinst4(
		.O(Q_out_dp4), // LUT general output
		.I0(Q_out_dp3) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_dpinst5(
		.O(Q_out_dp5), // LUT general output
		.I0(Q_out_dp4) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_dpinst6(
		.O(Q_out_dp6), // LUT general output
		.I0(Q_out_dp5) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_dpinst7(
		.O(Q_out_dp7), // LUT general output
		.I0(Q_out_dp6) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_dpinst8(
		.O(Q_out_dp8), // LUT general output
		.I0(Q_out_dp7) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_dpinst9(
		.O(Q_out_dp9), // LUT general output
		.I0(Q_out_dp8) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_dpinst10(
		.O(Q_out_dp10), // LUT general output
		.I0(Q_out_dp9) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_dpinst11(
		.O(Q_out_dp11), // LUT general output
		.I0(Q_out_dp10) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_dpinst12(
		.O(Q_out_dp12), // LUT general output
		.I0(Q_out_dp11) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_dpinst13(
		.O(Q_out_dp13), // LUT general output
		.I0(Q_out_dp12) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_dpinst14(
		.O(Q_out_dp14), // LUT general output
		.I0(Q_out_dp13) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_dpinst15(
		.O(Q_out_dp15), // LUT general output
		.I0(Q_out_dp14) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_dpinst16(
		.O(Q_out_dp16), // LUT general output
		.I0(Q_out_dp15) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_dpinst17(
		.O(Q_out_dp17), // LUT general output
		.I0(Q_out_dp16) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_dpinst18(
		.O(Q_out_dp18), // LUT general output
		.I0(Q_out_dp17) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_dpinst19(
		.O(Q_out_dp19), // LUT general output
		.I0(Q_out_dp18) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_dpinst20(
		.O(Q_out_dp20), // LUT general output
		.I0(Q_out_dp19) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_dpinst21(
		.O(Q_out_dp21), // LUT general output
		.I0(Q_out_dp20) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_dpinst22(
		.O(Q_out_dp22), // LUT general output
		.I0(Q_out_dp21) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_dpinst23(
		.O(Q_out_dp23), // LUT general output
		.I0(Q_out_dp22) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_dpinst24(
		.O(Q_out_dp24), // LUT general output
		.I0(Q_out_dp23) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_dpinst25(
		.O(Q_out_dp25), // LUT general output
		.I0(Q_out_dp24) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_dpinst26(
		.O(Q_out_dp26), // LUT general output
		.I0(Q_out_dp25) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_dpinst27(
		.O(Q_out_dp27), // LUT general output
		.I0(Q_out_dp26) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_dpinst28(
		.O(Q_out_dp28), // LUT general output
		.I0(Q_out_dp27) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_dpinst29(
		.O(Q_out_dp29), // LUT general output
		.I0(Q_out_dp28) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_dpinst30(
		.O(Q_out_dp30), // LUT general output
		.I0(Q_out_dp29) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_dpinst31(
		.O(Q_out_dp31), // LUT general output
		.I0(Q_out_dp30) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_dpinst32(
		.O(Q_out_dp32), // LUT general output
		.I0(Q_out_dp31) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_dpinst33(
		.O(Q_out_dp33), // LUT general output
		.I0(Q_out_dp32) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_dpinst34(
		.O(Q_out_dp34), // LUT general output
		.I0(Q_out_dp33) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_dpinst35(
		.O(Q_out_dp35), // LUT general output
		.I0(Q_out_dp34) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_dpinst36(
		.O(Q_out_dp36), // LUT general output
		.I0(Q_out_dp35) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_dpinst37(
		.O(Q_out_dp37), // LUT general output
		.I0(Q_out_dp36) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_dpinst38(
		.O(Q_out_dp38), // LUT general output
		.I0(Q_out_dp37) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_dpinst39(
		.O(Q_out_dp39), // LUT general output
		.I0(Q_out_dp38) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_dpinst40(
		.O(Q_out_dp40), // LUT general output
		.I0(Q_out_dp39) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_dpinst41(
		.O(Q_out_dp41), // LUT general output
		.I0(Q_out_dp40) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_dpinst42(
		.O(Q_out_dp42), // LUT general output
		.I0(Q_out_dp41) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_dpinst43(
		.O(Q_out_dp43), // LUT general output
		.I0(Q_out_dp42) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_dpinst44(
		.O(Q_out_dp44), // LUT general output
		.I0(Q_out_dp43) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_dpinst45(
		.O(Q_out_dp45), // LUT general output
		.I0(Q_out_dp44) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_dpinst46(
		.O(Q_out_dp46), // LUT general output
		.I0(Q_out_dp45) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_dpinst47(
		.O(Q_out_dp47), // LUT general output
		.I0(Q_out_dp46) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_dpinst48(
		.O(Q_out_dp48), // LUT general output
		.I0(Q_out_dp47) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_dpinst49(
		.O(Q_out_dp49), // LUT general output
		.I0(Q_out_dp48) // LUT input
	);

LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_dpinst50(
		.O(Q_out_dp50), // LUT general output
		.I0(Q_out_dp49) // LUT input
	);


LUT1 #(
		.INIT(2'b10) // Specify LUT Contents
		) LUT1_dpinst51(
		.O(delayed_edge), // LUT general output
		.I0(Q_out_dp50) // LUT input
	);



   //------------------------------------------------
   assign gpio_startn = ~blk_drdy;
   assign gpio_endn   = 1'b0; //~blk_dvld;
   assign gpio_exec   = 1'b0; //blk_busy;
	

   always @(posedge clk) blk_drdy_delay <= blk_drdy;

   AES_Composite_enc AES_Composite_enc
     (.Kin(blk_kin), .Din(blk_din), .Dout(blk_dout),
      .Krdy(blk_krdy), .Drdy(blk_drdy_delay), .Kvld(blk_kvld), .Dvld(blk_dvld),
      /*.EncDec(blk_encdec),*/ .EN(blk_en), .BSY(blk_busy),
		.CLK_IN(Q_out3), .RSTn(blk_rstn), .stop_detect(stop_detect), .delayed_edge(delayed_edge));

// BT: 	Q_out3 is the intended slightly delayed clock for our AES system
//			it is the output of 'clk_delay' in paper (Figure 4)

   //------------------------------------------------   
   MK_CLKRST mk_clkrst (.clkin(lbus_clkn), .rstnin(lbus_rstn),
                        .clk(clk), .rst(rst));
endmodule // CHIP_SASEBO_GIII_AES


   
//================================================ MK_CLKRST
module MK_CLKRST (clkin, rstnin, clk, rst);
   //synthesis attribute keep_hierarchy of MK_CLKRST is no;
   
   //------------------------------------------------
   input  clkin, rstnin;
   output clk, rst;
   
   //------------------------------------------------
   wire   refclk;
//   wire   clk_dcm, locked;

   //------------------------------------------------ clock
   IBUFG u10 (.I(clkin), .O(refclk)); 
   BUFG  u12 (.I(refclk),   .O(clk));

   //------------------------------------------------ reset
   MK_RST u20 (.locked(rstnin), .clk(clk), .rst(rst));
endmodule // MK_CLKRST



//================================================ MK_RST
module MK_RST (locked, clk, rst);
   //synthesis attribute keep_hierarchy of MK_RST is no;
   
   //------------------------------------------------
   input  locked, clk;
   output rst;

   //------------------------------------------------
   reg [15:0] cnt;
   
   //------------------------------------------------
   always @(posedge clk or negedge locked) 
     if (~locked)    cnt <= 16'h0;
     else if (~&cnt) cnt <= cnt + 16'h1;

   assign rst = ~&cnt;
endmodule // MK_RST
